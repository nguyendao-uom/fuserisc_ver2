	//External IO ports exported directly from the corresponding tiles
module eFPGA (Tile_X4Y1_OPA_I0, Tile_X4Y1_OPA_I1, Tile_X4Y1_OPA_I2, Tile_X4Y1_OPA_I3, UserCLK, Tile_X4Y1_OPB_I0, Tile_X4Y1_OPB_I1, Tile_X4Y1_OPB_I2, Tile_X4Y1_OPB_I3, Tile_X4Y1_RES0_O0, Tile_X4Y1_RES0_O1, Tile_X4Y1_RES0_O2, Tile_X4Y1_RES0_O3, Tile_X4Y1_RES1_O0, Tile_X4Y1_RES1_O1, Tile_X4Y1_RES1_O2, Tile_X4Y1_RES1_O3, Tile_X4Y1_RES2_O0, Tile_X4Y1_RES2_O1, Tile_X4Y1_RES2_O2, Tile_X4Y1_RES2_O3, Tile_X11Y1_OPA_I0, Tile_X11Y1_OPA_I1, Tile_X11Y1_OPA_I2, Tile_X11Y1_OPA_I3, Tile_X11Y1_OPB_I0, Tile_X11Y1_OPB_I1, Tile_X11Y1_OPB_I2, Tile_X11Y1_OPB_I3, Tile_X11Y1_RES0_O0, Tile_X11Y1_RES0_O1, Tile_X11Y1_RES0_O2, Tile_X11Y1_RES0_O3, Tile_X11Y1_RES1_O0, Tile_X11Y1_RES1_O1, Tile_X11Y1_RES1_O2, Tile_X11Y1_RES1_O3, Tile_X11Y1_RES2_O0, Tile_X11Y1_RES2_O1, Tile_X11Y1_RES2_O2, Tile_X11Y1_RES2_O3, Tile_X4Y2_OPA_I0, Tile_X4Y2_OPA_I1, Tile_X4Y2_OPA_I2, Tile_X4Y2_OPA_I3, Tile_X4Y2_OPB_I0, Tile_X4Y2_OPB_I1, Tile_X4Y2_OPB_I2, Tile_X4Y2_OPB_I3, Tile_X4Y2_RES0_O0, Tile_X4Y2_RES0_O1, Tile_X4Y2_RES0_O2, Tile_X4Y2_RES0_O3, Tile_X4Y2_RES1_O0, Tile_X4Y2_RES1_O1, Tile_X4Y2_RES1_O2, Tile_X4Y2_RES1_O3, Tile_X4Y2_RES2_O0, Tile_X4Y2_RES2_O1, Tile_X4Y2_RES2_O2, Tile_X4Y2_RES2_O3, Tile_X11Y2_OPA_I0, Tile_X11Y2_OPA_I1, Tile_X11Y2_OPA_I2, Tile_X11Y2_OPA_I3, Tile_X11Y2_OPB_I0, Tile_X11Y2_OPB_I1, Tile_X11Y2_OPB_I2, Tile_X11Y2_OPB_I3, Tile_X11Y2_RES0_O0, Tile_X11Y2_RES0_O1, Tile_X11Y2_RES0_O2, Tile_X11Y2_RES0_O3, Tile_X11Y2_RES1_O0, Tile_X11Y2_RES1_O1, Tile_X11Y2_RES1_O2, Tile_X11Y2_RES1_O3, Tile_X11Y2_RES2_O0, Tile_X11Y2_RES2_O1, Tile_X11Y2_RES2_O2, Tile_X11Y2_RES2_O3, Tile_X4Y3_OPA_I0, Tile_X4Y3_OPA_I1, Tile_X4Y3_OPA_I2, Tile_X4Y3_OPA_I3, Tile_X4Y3_OPB_I0, Tile_X4Y3_OPB_I1, Tile_X4Y3_OPB_I2, Tile_X4Y3_OPB_I3, Tile_X4Y3_RES0_O0, Tile_X4Y3_RES0_O1, Tile_X4Y3_RES0_O2, Tile_X4Y3_RES0_O3, Tile_X4Y3_RES1_O0, Tile_X4Y3_RES1_O1, Tile_X4Y3_RES1_O2, Tile_X4Y3_RES1_O3, Tile_X4Y3_RES2_O0, Tile_X4Y3_RES2_O1, Tile_X4Y3_RES2_O2, Tile_X4Y3_RES2_O3, Tile_X11Y3_OPA_I0, Tile_X11Y3_OPA_I1, Tile_X11Y3_OPA_I2, Tile_X11Y3_OPA_I3, Tile_X11Y3_OPB_I0, Tile_X11Y3_OPB_I1, Tile_X11Y3_OPB_I2, Tile_X11Y3_OPB_I3, Tile_X11Y3_RES0_O0, Tile_X11Y3_RES0_O1, Tile_X11Y3_RES0_O2, Tile_X11Y3_RES0_O3, Tile_X11Y3_RES1_O0, Tile_X11Y3_RES1_O1, Tile_X11Y3_RES1_O2, Tile_X11Y3_RES1_O3, Tile_X11Y3_RES2_O0, Tile_X11Y3_RES2_O1, Tile_X11Y3_RES2_O2, Tile_X11Y3_RES2_O3, Tile_X4Y4_OPA_I0, Tile_X4Y4_OPA_I1, Tile_X4Y4_OPA_I2, Tile_X4Y4_OPA_I3, Tile_X4Y4_OPB_I0, Tile_X4Y4_OPB_I1, Tile_X4Y4_OPB_I2, Tile_X4Y4_OPB_I3, Tile_X4Y4_RES0_O0, Tile_X4Y4_RES0_O1, Tile_X4Y4_RES0_O2, Tile_X4Y4_RES0_O3, Tile_X4Y4_RES1_O0, Tile_X4Y4_RES1_O1, Tile_X4Y4_RES1_O2, Tile_X4Y4_RES1_O3, Tile_X4Y4_RES2_O0, Tile_X4Y4_RES2_O1, Tile_X4Y4_RES2_O2, Tile_X4Y4_RES2_O3, Tile_X11Y4_OPA_I0, Tile_X11Y4_OPA_I1, Tile_X11Y4_OPA_I2, Tile_X11Y4_OPA_I3, Tile_X11Y4_OPB_I0, Tile_X11Y4_OPB_I1, Tile_X11Y4_OPB_I2, Tile_X11Y4_OPB_I3, Tile_X11Y4_RES0_O0, Tile_X11Y4_RES0_O1, Tile_X11Y4_RES0_O2, Tile_X11Y4_RES0_O3, Tile_X11Y4_RES1_O0, Tile_X11Y4_RES1_O1, Tile_X11Y4_RES1_O2, Tile_X11Y4_RES1_O3, Tile_X11Y4_RES2_O0, Tile_X11Y4_RES2_O1, Tile_X11Y4_RES2_O2, Tile_X11Y4_RES2_O3, Tile_X4Y5_OPA_I0, Tile_X4Y5_OPA_I1, Tile_X4Y5_OPA_I2, Tile_X4Y5_OPA_I3, Tile_X4Y5_OPB_I0, Tile_X4Y5_OPB_I1, Tile_X4Y5_OPB_I2, Tile_X4Y5_OPB_I3, Tile_X4Y5_RES0_O0, Tile_X4Y5_RES0_O1, Tile_X4Y5_RES0_O2, Tile_X4Y5_RES0_O3, Tile_X4Y5_RES1_O0, Tile_X4Y5_RES1_O1, Tile_X4Y5_RES1_O2, Tile_X4Y5_RES1_O3, Tile_X4Y5_RES2_O0, Tile_X4Y5_RES2_O1, Tile_X4Y5_RES2_O2, Tile_X4Y5_RES2_O3, Tile_X11Y5_OPA_I0, Tile_X11Y5_OPA_I1, Tile_X11Y5_OPA_I2, Tile_X11Y5_OPA_I3, Tile_X11Y5_OPB_I0, Tile_X11Y5_OPB_I1, Tile_X11Y5_OPB_I2, Tile_X11Y5_OPB_I3, Tile_X11Y5_RES0_O0, Tile_X11Y5_RES0_O1, Tile_X11Y5_RES0_O2, Tile_X11Y5_RES0_O3, Tile_X11Y5_RES1_O0, Tile_X11Y5_RES1_O1, Tile_X11Y5_RES1_O2, Tile_X11Y5_RES1_O3, Tile_X11Y5_RES2_O0, Tile_X11Y5_RES2_O1, Tile_X11Y5_RES2_O2, Tile_X11Y5_RES2_O3, Tile_X4Y6_OPA_I0, Tile_X4Y6_OPA_I1, Tile_X4Y6_OPA_I2, Tile_X4Y6_OPA_I3, Tile_X4Y6_OPB_I0, Tile_X4Y6_OPB_I1, Tile_X4Y6_OPB_I2, Tile_X4Y6_OPB_I3, Tile_X4Y6_RES0_O0, Tile_X4Y6_RES0_O1, Tile_X4Y6_RES0_O2, Tile_X4Y6_RES0_O3, Tile_X4Y6_RES1_O0, Tile_X4Y6_RES1_O1, Tile_X4Y6_RES1_O2, Tile_X4Y6_RES1_O3, Tile_X4Y6_RES2_O0, Tile_X4Y6_RES2_O1, Tile_X4Y6_RES2_O2, Tile_X4Y6_RES2_O3, Tile_X11Y6_OPA_I0, Tile_X11Y6_OPA_I1, Tile_X11Y6_OPA_I2, Tile_X11Y6_OPA_I3, Tile_X11Y6_OPB_I0, Tile_X11Y6_OPB_I1, Tile_X11Y6_OPB_I2, Tile_X11Y6_OPB_I3, Tile_X11Y6_RES0_O0, Tile_X11Y6_RES0_O1, Tile_X11Y6_RES0_O2, Tile_X11Y6_RES0_O3, Tile_X11Y6_RES1_O0, Tile_X11Y6_RES1_O1, Tile_X11Y6_RES1_O2, Tile_X11Y6_RES1_O3, Tile_X11Y6_RES2_O0, Tile_X11Y6_RES2_O1, Tile_X11Y6_RES2_O2, Tile_X11Y6_RES2_O3, Tile_X4Y7_OPA_I0, Tile_X4Y7_OPA_I1, Tile_X4Y7_OPA_I2, Tile_X4Y7_OPA_I3, Tile_X4Y7_OPB_I0, Tile_X4Y7_OPB_I1, Tile_X4Y7_OPB_I2, Tile_X4Y7_OPB_I3, Tile_X4Y7_RES0_O0, Tile_X4Y7_RES0_O1, Tile_X4Y7_RES0_O2, Tile_X4Y7_RES0_O3, Tile_X4Y7_RES1_O0, Tile_X4Y7_RES1_O1, Tile_X4Y7_RES1_O2, Tile_X4Y7_RES1_O3, Tile_X4Y7_RES2_O0, Tile_X4Y7_RES2_O1, Tile_X4Y7_RES2_O2, Tile_X4Y7_RES2_O3, Tile_X11Y7_OPA_I0, Tile_X11Y7_OPA_I1, Tile_X11Y7_OPA_I2, Tile_X11Y7_OPA_I3, Tile_X11Y7_OPB_I0, Tile_X11Y7_OPB_I1, Tile_X11Y7_OPB_I2, Tile_X11Y7_OPB_I3, Tile_X11Y7_RES0_O0, Tile_X11Y7_RES0_O1, Tile_X11Y7_RES0_O2, Tile_X11Y7_RES0_O3, Tile_X11Y7_RES1_O0, Tile_X11Y7_RES1_O1, Tile_X11Y7_RES1_O2, Tile_X11Y7_RES1_O3, Tile_X11Y7_RES2_O0, Tile_X11Y7_RES2_O1, Tile_X11Y7_RES2_O2, Tile_X11Y7_RES2_O3, Tile_X4Y8_OPA_I0, Tile_X4Y8_OPA_I1, Tile_X4Y8_OPA_I2, Tile_X4Y8_OPA_I3, Tile_X4Y8_OPB_I0, Tile_X4Y8_OPB_I1, Tile_X4Y8_OPB_I2, Tile_X4Y8_OPB_I3, Tile_X4Y8_RES0_O0, Tile_X4Y8_RES0_O1, Tile_X4Y8_RES0_O2, Tile_X4Y8_RES0_O3, Tile_X4Y8_RES1_O0, Tile_X4Y8_RES1_O1, Tile_X4Y8_RES1_O2, Tile_X4Y8_RES1_O3, Tile_X4Y8_RES2_O0, Tile_X4Y8_RES2_O1, Tile_X4Y8_RES2_O2, Tile_X4Y8_RES2_O3, Tile_X11Y8_OPA_I0, Tile_X11Y8_OPA_I1, Tile_X11Y8_OPA_I2, Tile_X11Y8_OPA_I3, Tile_X11Y8_OPB_I0, Tile_X11Y8_OPB_I1, Tile_X11Y8_OPB_I2, Tile_X11Y8_OPB_I3, Tile_X11Y8_RES0_O0, Tile_X11Y8_RES0_O1, Tile_X11Y8_RES0_O2, Tile_X11Y8_RES0_O3, Tile_X11Y8_RES1_O0, Tile_X11Y8_RES1_O1, Tile_X11Y8_RES1_O2, Tile_X11Y8_RES1_O3, Tile_X11Y8_RES2_O0, Tile_X11Y8_RES2_O1, Tile_X11Y8_RES2_O2, Tile_X11Y8_RES2_O3, Tile_X4Y9_OPA_I0, Tile_X4Y9_OPA_I1, Tile_X4Y9_OPA_I2, Tile_X4Y9_OPA_I3, Tile_X4Y9_OPB_I0, Tile_X4Y9_OPB_I1, Tile_X4Y9_OPB_I2, Tile_X4Y9_OPB_I3, Tile_X4Y9_RES0_O0, Tile_X4Y9_RES0_O1, Tile_X4Y9_RES0_O2, Tile_X4Y9_RES0_O3, Tile_X4Y9_RES1_O0, Tile_X4Y9_RES1_O1, Tile_X4Y9_RES1_O2, Tile_X4Y9_RES1_O3, Tile_X4Y9_RES2_O0, Tile_X4Y9_RES2_O1, Tile_X4Y9_RES2_O2, Tile_X4Y9_RES2_O3, Tile_X11Y9_OPA_I0, Tile_X11Y9_OPA_I1, Tile_X11Y9_OPA_I2, Tile_X11Y9_OPA_I3, Tile_X11Y9_OPB_I0, Tile_X11Y9_OPB_I1, Tile_X11Y9_OPB_I2, Tile_X11Y9_OPB_I3, Tile_X11Y9_RES0_O0, Tile_X11Y9_RES0_O1, Tile_X11Y9_RES0_O2, Tile_X11Y9_RES0_O3, Tile_X11Y9_RES1_O0, Tile_X11Y9_RES1_O1, Tile_X11Y9_RES1_O2, Tile_X11Y9_RES1_O3, Tile_X11Y9_RES2_O0, Tile_X11Y9_RES2_O1, Tile_X11Y9_RES2_O2, Tile_X11Y9_RES2_O3, Tile_X0Y10_A_I_top, Tile_X0Y10_A_T_top, Tile_X0Y10_A_O_top, Tile_X0Y10_B_I_top, Tile_X0Y10_B_T_top, Tile_X0Y10_B_O_top, Tile_X0Y10_A_config_C_bit0, Tile_X0Y10_A_config_C_bit1, Tile_X0Y10_A_config_C_bit2, Tile_X0Y10_A_config_C_bit3, Tile_X0Y10_B_config_C_bit0, Tile_X0Y10_B_config_C_bit1, Tile_X0Y10_B_config_C_bit2, Tile_X0Y10_B_config_C_bit3, Tile_X15Y10_RAM2FAB_D0_I0, Tile_X15Y10_RAM2FAB_D0_I1, Tile_X15Y10_RAM2FAB_D0_I2, Tile_X15Y10_RAM2FAB_D0_I3, Tile_X15Y10_RAM2FAB_D1_I0, Tile_X15Y10_RAM2FAB_D1_I1, Tile_X15Y10_RAM2FAB_D1_I2, Tile_X15Y10_RAM2FAB_D1_I3, Tile_X15Y10_RAM2FAB_D2_I0, Tile_X15Y10_RAM2FAB_D2_I1, Tile_X15Y10_RAM2FAB_D2_I2, Tile_X15Y10_RAM2FAB_D2_I3, Tile_X15Y10_RAM2FAB_D3_I0, Tile_X15Y10_RAM2FAB_D3_I1, Tile_X15Y10_RAM2FAB_D3_I2, Tile_X15Y10_RAM2FAB_D3_I3, Tile_X15Y10_FAB2RAM_D0_O0, Tile_X15Y10_FAB2RAM_D0_O1, Tile_X15Y10_FAB2RAM_D0_O2, Tile_X15Y10_FAB2RAM_D0_O3, Tile_X15Y10_FAB2RAM_D1_O0, Tile_X15Y10_FAB2RAM_D1_O1, Tile_X15Y10_FAB2RAM_D1_O2, Tile_X15Y10_FAB2RAM_D1_O3, Tile_X15Y10_FAB2RAM_D2_O0, Tile_X15Y10_FAB2RAM_D2_O1, Tile_X15Y10_FAB2RAM_D2_O2, Tile_X15Y10_FAB2RAM_D2_O3, Tile_X15Y10_FAB2RAM_D3_O0, Tile_X15Y10_FAB2RAM_D3_O1, Tile_X15Y10_FAB2RAM_D3_O2, Tile_X15Y10_FAB2RAM_D3_O3, Tile_X15Y10_FAB2RAM_A0_O0, Tile_X15Y10_FAB2RAM_A0_O1, Tile_X15Y10_FAB2RAM_A0_O2, Tile_X15Y10_FAB2RAM_A0_O3, Tile_X15Y10_FAB2RAM_A1_O0, Tile_X15Y10_FAB2RAM_A1_O1, Tile_X15Y10_FAB2RAM_A1_O2, Tile_X15Y10_FAB2RAM_A1_O3, Tile_X15Y10_FAB2RAM_C_O0, Tile_X15Y10_FAB2RAM_C_O1, Tile_X15Y10_FAB2RAM_C_O2, Tile_X15Y10_FAB2RAM_C_O3, Tile_X15Y10_Config_accessC_bit0, Tile_X15Y10_Config_accessC_bit1, Tile_X15Y10_Config_accessC_bit2, Tile_X15Y10_Config_accessC_bit3, Tile_X0Y11_A_I_top, Tile_X0Y11_A_T_top, Tile_X0Y11_A_O_top, Tile_X0Y11_B_I_top, Tile_X0Y11_B_T_top, Tile_X0Y11_B_O_top, Tile_X0Y11_A_config_C_bit0, Tile_X0Y11_A_config_C_bit1, Tile_X0Y11_A_config_C_bit2, Tile_X0Y11_A_config_C_bit3, Tile_X0Y11_B_config_C_bit0, Tile_X0Y11_B_config_C_bit1, Tile_X0Y11_B_config_C_bit2, Tile_X0Y11_B_config_C_bit3, Tile_X15Y11_RAM2FAB_D0_I0, Tile_X15Y11_RAM2FAB_D0_I1, Tile_X15Y11_RAM2FAB_D0_I2, Tile_X15Y11_RAM2FAB_D0_I3, Tile_X15Y11_RAM2FAB_D1_I0, Tile_X15Y11_RAM2FAB_D1_I1, Tile_X15Y11_RAM2FAB_D1_I2, Tile_X15Y11_RAM2FAB_D1_I3, Tile_X15Y11_RAM2FAB_D2_I0, Tile_X15Y11_RAM2FAB_D2_I1, Tile_X15Y11_RAM2FAB_D2_I2, Tile_X15Y11_RAM2FAB_D2_I3, Tile_X15Y11_RAM2FAB_D3_I0, Tile_X15Y11_RAM2FAB_D3_I1, Tile_X15Y11_RAM2FAB_D3_I2, Tile_X15Y11_RAM2FAB_D3_I3, Tile_X15Y11_FAB2RAM_D0_O0, Tile_X15Y11_FAB2RAM_D0_O1, Tile_X15Y11_FAB2RAM_D0_O2, Tile_X15Y11_FAB2RAM_D0_O3, Tile_X15Y11_FAB2RAM_D1_O0, Tile_X15Y11_FAB2RAM_D1_O1, Tile_X15Y11_FAB2RAM_D1_O2, Tile_X15Y11_FAB2RAM_D1_O3, Tile_X15Y11_FAB2RAM_D2_O0, Tile_X15Y11_FAB2RAM_D2_O1, Tile_X15Y11_FAB2RAM_D2_O2, Tile_X15Y11_FAB2RAM_D2_O3, Tile_X15Y11_FAB2RAM_D3_O0, Tile_X15Y11_FAB2RAM_D3_O1, Tile_X15Y11_FAB2RAM_D3_O2, Tile_X15Y11_FAB2RAM_D3_O3, Tile_X15Y11_FAB2RAM_A0_O0, Tile_X15Y11_FAB2RAM_A0_O1, Tile_X15Y11_FAB2RAM_A0_O2, Tile_X15Y11_FAB2RAM_A0_O3, Tile_X15Y11_FAB2RAM_A1_O0, Tile_X15Y11_FAB2RAM_A1_O1, Tile_X15Y11_FAB2RAM_A1_O2, Tile_X15Y11_FAB2RAM_A1_O3, Tile_X15Y11_FAB2RAM_C_O0, Tile_X15Y11_FAB2RAM_C_O1, Tile_X15Y11_FAB2RAM_C_O2, Tile_X15Y11_FAB2RAM_C_O3, Tile_X15Y11_Config_accessC_bit0, Tile_X15Y11_Config_accessC_bit1, Tile_X15Y11_Config_accessC_bit2, Tile_X15Y11_Config_accessC_bit3, Tile_X0Y12_A_I_top, Tile_X0Y12_A_T_top, Tile_X0Y12_A_O_top, Tile_X0Y12_B_I_top, Tile_X0Y12_B_T_top, Tile_X0Y12_B_O_top, Tile_X0Y12_A_config_C_bit0, Tile_X0Y12_A_config_C_bit1, Tile_X0Y12_A_config_C_bit2, Tile_X0Y12_A_config_C_bit3, Tile_X0Y12_B_config_C_bit0, Tile_X0Y12_B_config_C_bit1, Tile_X0Y12_B_config_C_bit2, Tile_X0Y12_B_config_C_bit3, Tile_X15Y12_RAM2FAB_D0_I0, Tile_X15Y12_RAM2FAB_D0_I1, Tile_X15Y12_RAM2FAB_D0_I2, Tile_X15Y12_RAM2FAB_D0_I3, Tile_X15Y12_RAM2FAB_D1_I0, Tile_X15Y12_RAM2FAB_D1_I1, Tile_X15Y12_RAM2FAB_D1_I2, Tile_X15Y12_RAM2FAB_D1_I3, Tile_X15Y12_RAM2FAB_D2_I0, Tile_X15Y12_RAM2FAB_D2_I1, Tile_X15Y12_RAM2FAB_D2_I2, Tile_X15Y12_RAM2FAB_D2_I3, Tile_X15Y12_RAM2FAB_D3_I0, Tile_X15Y12_RAM2FAB_D3_I1, Tile_X15Y12_RAM2FAB_D3_I2, Tile_X15Y12_RAM2FAB_D3_I3, Tile_X15Y12_FAB2RAM_D0_O0, Tile_X15Y12_FAB2RAM_D0_O1, Tile_X15Y12_FAB2RAM_D0_O2, Tile_X15Y12_FAB2RAM_D0_O3, Tile_X15Y12_FAB2RAM_D1_O0, Tile_X15Y12_FAB2RAM_D1_O1, Tile_X15Y12_FAB2RAM_D1_O2, Tile_X15Y12_FAB2RAM_D1_O3, Tile_X15Y12_FAB2RAM_D2_O0, Tile_X15Y12_FAB2RAM_D2_O1, Tile_X15Y12_FAB2RAM_D2_O2, Tile_X15Y12_FAB2RAM_D2_O3, Tile_X15Y12_FAB2RAM_D3_O0, Tile_X15Y12_FAB2RAM_D3_O1, Tile_X15Y12_FAB2RAM_D3_O2, Tile_X15Y12_FAB2RAM_D3_O3, Tile_X15Y12_FAB2RAM_A0_O0, Tile_X15Y12_FAB2RAM_A0_O1, Tile_X15Y12_FAB2RAM_A0_O2, Tile_X15Y12_FAB2RAM_A0_O3, Tile_X15Y12_FAB2RAM_A1_O0, Tile_X15Y12_FAB2RAM_A1_O1, Tile_X15Y12_FAB2RAM_A1_O2, Tile_X15Y12_FAB2RAM_A1_O3, Tile_X15Y12_FAB2RAM_C_O0, Tile_X15Y12_FAB2RAM_C_O1, Tile_X15Y12_FAB2RAM_C_O2, Tile_X15Y12_FAB2RAM_C_O3, Tile_X15Y12_Config_accessC_bit0, Tile_X15Y12_Config_accessC_bit1, Tile_X15Y12_Config_accessC_bit2, Tile_X15Y12_Config_accessC_bit3, FrameData, FrameStrobe);
	parameter MaxFramesPerCol = 20;
	parameter FrameBitsPerRow = 32;
	parameter NoConfigBits = 0;
	input Tile_X4Y1_OPA_I0;  //EXTERNAL
	input Tile_X4Y1_OPA_I1;  //EXTERNAL
	input Tile_X4Y1_OPA_I2;  //EXTERNAL
	input Tile_X4Y1_OPA_I3;  //EXTERNAL
	input UserCLK;  //EXTERNAL //SHARED_PORT //## the EXTERNAL keyword will send this signal all the way to top and the --SHARED Allows multiple BELs usg the same port (e.g. for exportg a clock to the top)
	input Tile_X4Y1_OPB_I0;  //EXTERNAL
	input Tile_X4Y1_OPB_I1;  //EXTERNAL
	input Tile_X4Y1_OPB_I2;  //EXTERNAL
	input Tile_X4Y1_OPB_I3;  //EXTERNAL
	output Tile_X4Y1_RES0_O0;  //EXTERNAL
	output Tile_X4Y1_RES0_O1;  //EXTERNAL
	output Tile_X4Y1_RES0_O2;  //EXTERNAL
	output Tile_X4Y1_RES0_O3;  //EXTERNAL
	output Tile_X4Y1_RES1_O0;  //EXTERNAL
	output Tile_X4Y1_RES1_O1;  //EXTERNAL
	output Tile_X4Y1_RES1_O2;  //EXTERNAL
	output Tile_X4Y1_RES1_O3;  //EXTERNAL
	output Tile_X4Y1_RES2_O0;  //EXTERNAL
	output Tile_X4Y1_RES2_O1;  //EXTERNAL
	output Tile_X4Y1_RES2_O2;  //EXTERNAL
	output Tile_X4Y1_RES2_O3;  //EXTERNAL
	input Tile_X11Y1_OPA_I0;  //EXTERNAL
	input Tile_X11Y1_OPA_I1;  //EXTERNAL
	input Tile_X11Y1_OPA_I2;  //EXTERNAL
	input Tile_X11Y1_OPA_I3;  //EXTERNAL
	input Tile_X11Y1_OPB_I0;  //EXTERNAL
	input Tile_X11Y1_OPB_I1;  //EXTERNAL
	input Tile_X11Y1_OPB_I2;  //EXTERNAL
	input Tile_X11Y1_OPB_I3;  //EXTERNAL
	output Tile_X11Y1_RES0_O0;  //EXTERNAL
	output Tile_X11Y1_RES0_O1;  //EXTERNAL
	output Tile_X11Y1_RES0_O2;  //EXTERNAL
	output Tile_X11Y1_RES0_O3;  //EXTERNAL
	output Tile_X11Y1_RES1_O0;  //EXTERNAL
	output Tile_X11Y1_RES1_O1;  //EXTERNAL
	output Tile_X11Y1_RES1_O2;  //EXTERNAL
	output Tile_X11Y1_RES1_O3;  //EXTERNAL
	output Tile_X11Y1_RES2_O0;  //EXTERNAL
	output Tile_X11Y1_RES2_O1;  //EXTERNAL
	output Tile_X11Y1_RES2_O2;  //EXTERNAL
	output Tile_X11Y1_RES2_O3;  //EXTERNAL
	input Tile_X4Y2_OPA_I0;  //EXTERNAL
	input Tile_X4Y2_OPA_I1;  //EXTERNAL
	input Tile_X4Y2_OPA_I2;  //EXTERNAL
	input Tile_X4Y2_OPA_I3;  //EXTERNAL
	input Tile_X4Y2_OPB_I0;  //EXTERNAL
	input Tile_X4Y2_OPB_I1;  //EXTERNAL
	input Tile_X4Y2_OPB_I2;  //EXTERNAL
	input Tile_X4Y2_OPB_I3;  //EXTERNAL
	output Tile_X4Y2_RES0_O0;  //EXTERNAL
	output Tile_X4Y2_RES0_O1;  //EXTERNAL
	output Tile_X4Y2_RES0_O2;  //EXTERNAL
	output Tile_X4Y2_RES0_O3;  //EXTERNAL
	output Tile_X4Y2_RES1_O0;  //EXTERNAL
	output Tile_X4Y2_RES1_O1;  //EXTERNAL
	output Tile_X4Y2_RES1_O2;  //EXTERNAL
	output Tile_X4Y2_RES1_O3;  //EXTERNAL
	output Tile_X4Y2_RES2_O0;  //EXTERNAL
	output Tile_X4Y2_RES2_O1;  //EXTERNAL
	output Tile_X4Y2_RES2_O2;  //EXTERNAL
	output Tile_X4Y2_RES2_O3;  //EXTERNAL
	input Tile_X11Y2_OPA_I0;  //EXTERNAL
	input Tile_X11Y2_OPA_I1;  //EXTERNAL
	input Tile_X11Y2_OPA_I2;  //EXTERNAL
	input Tile_X11Y2_OPA_I3;  //EXTERNAL
	input Tile_X11Y2_OPB_I0;  //EXTERNAL
	input Tile_X11Y2_OPB_I1;  //EXTERNAL
	input Tile_X11Y2_OPB_I2;  //EXTERNAL
	input Tile_X11Y2_OPB_I3;  //EXTERNAL
	output Tile_X11Y2_RES0_O0;  //EXTERNAL
	output Tile_X11Y2_RES0_O1;  //EXTERNAL
	output Tile_X11Y2_RES0_O2;  //EXTERNAL
	output Tile_X11Y2_RES0_O3;  //EXTERNAL
	output Tile_X11Y2_RES1_O0;  //EXTERNAL
	output Tile_X11Y2_RES1_O1;  //EXTERNAL
	output Tile_X11Y2_RES1_O2;  //EXTERNAL
	output Tile_X11Y2_RES1_O3;  //EXTERNAL
	output Tile_X11Y2_RES2_O0;  //EXTERNAL
	output Tile_X11Y2_RES2_O1;  //EXTERNAL
	output Tile_X11Y2_RES2_O2;  //EXTERNAL
	output Tile_X11Y2_RES2_O3;  //EXTERNAL
	input Tile_X4Y3_OPA_I0;  //EXTERNAL
	input Tile_X4Y3_OPA_I1;  //EXTERNAL
	input Tile_X4Y3_OPA_I2;  //EXTERNAL
	input Tile_X4Y3_OPA_I3;  //EXTERNAL
	input Tile_X4Y3_OPB_I0;  //EXTERNAL
	input Tile_X4Y3_OPB_I1;  //EXTERNAL
	input Tile_X4Y3_OPB_I2;  //EXTERNAL
	input Tile_X4Y3_OPB_I3;  //EXTERNAL
	output Tile_X4Y3_RES0_O0;  //EXTERNAL
	output Tile_X4Y3_RES0_O1;  //EXTERNAL
	output Tile_X4Y3_RES0_O2;  //EXTERNAL
	output Tile_X4Y3_RES0_O3;  //EXTERNAL
	output Tile_X4Y3_RES1_O0;  //EXTERNAL
	output Tile_X4Y3_RES1_O1;  //EXTERNAL
	output Tile_X4Y3_RES1_O2;  //EXTERNAL
	output Tile_X4Y3_RES1_O3;  //EXTERNAL
	output Tile_X4Y3_RES2_O0;  //EXTERNAL
	output Tile_X4Y3_RES2_O1;  //EXTERNAL
	output Tile_X4Y3_RES2_O2;  //EXTERNAL
	output Tile_X4Y3_RES2_O3;  //EXTERNAL
	input Tile_X11Y3_OPA_I0;  //EXTERNAL
	input Tile_X11Y3_OPA_I1;  //EXTERNAL
	input Tile_X11Y3_OPA_I2;  //EXTERNAL
	input Tile_X11Y3_OPA_I3;  //EXTERNAL
	input Tile_X11Y3_OPB_I0;  //EXTERNAL
	input Tile_X11Y3_OPB_I1;  //EXTERNAL
	input Tile_X11Y3_OPB_I2;  //EXTERNAL
	input Tile_X11Y3_OPB_I3;  //EXTERNAL
	output Tile_X11Y3_RES0_O0;  //EXTERNAL
	output Tile_X11Y3_RES0_O1;  //EXTERNAL
	output Tile_X11Y3_RES0_O2;  //EXTERNAL
	output Tile_X11Y3_RES0_O3;  //EXTERNAL
	output Tile_X11Y3_RES1_O0;  //EXTERNAL
	output Tile_X11Y3_RES1_O1;  //EXTERNAL
	output Tile_X11Y3_RES1_O2;  //EXTERNAL
	output Tile_X11Y3_RES1_O3;  //EXTERNAL
	output Tile_X11Y3_RES2_O0;  //EXTERNAL
	output Tile_X11Y3_RES2_O1;  //EXTERNAL
	output Tile_X11Y3_RES2_O2;  //EXTERNAL
	output Tile_X11Y3_RES2_O3;  //EXTERNAL
	input Tile_X4Y4_OPA_I0;  //EXTERNAL
	input Tile_X4Y4_OPA_I1;  //EXTERNAL
	input Tile_X4Y4_OPA_I2;  //EXTERNAL
	input Tile_X4Y4_OPA_I3;  //EXTERNAL
	input Tile_X4Y4_OPB_I0;  //EXTERNAL
	input Tile_X4Y4_OPB_I1;  //EXTERNAL
	input Tile_X4Y4_OPB_I2;  //EXTERNAL
	input Tile_X4Y4_OPB_I3;  //EXTERNAL
	output Tile_X4Y4_RES0_O0;  //EXTERNAL
	output Tile_X4Y4_RES0_O1;  //EXTERNAL
	output Tile_X4Y4_RES0_O2;  //EXTERNAL
	output Tile_X4Y4_RES0_O3;  //EXTERNAL
	output Tile_X4Y4_RES1_O0;  //EXTERNAL
	output Tile_X4Y4_RES1_O1;  //EXTERNAL
	output Tile_X4Y4_RES1_O2;  //EXTERNAL
	output Tile_X4Y4_RES1_O3;  //EXTERNAL
	output Tile_X4Y4_RES2_O0;  //EXTERNAL
	output Tile_X4Y4_RES2_O1;  //EXTERNAL
	output Tile_X4Y4_RES2_O2;  //EXTERNAL
	output Tile_X4Y4_RES2_O3;  //EXTERNAL
	input Tile_X11Y4_OPA_I0;  //EXTERNAL
	input Tile_X11Y4_OPA_I1;  //EXTERNAL
	input Tile_X11Y4_OPA_I2;  //EXTERNAL
	input Tile_X11Y4_OPA_I3;  //EXTERNAL
	input Tile_X11Y4_OPB_I0;  //EXTERNAL
	input Tile_X11Y4_OPB_I1;  //EXTERNAL
	input Tile_X11Y4_OPB_I2;  //EXTERNAL
	input Tile_X11Y4_OPB_I3;  //EXTERNAL
	output Tile_X11Y4_RES0_O0;  //EXTERNAL
	output Tile_X11Y4_RES0_O1;  //EXTERNAL
	output Tile_X11Y4_RES0_O2;  //EXTERNAL
	output Tile_X11Y4_RES0_O3;  //EXTERNAL
	output Tile_X11Y4_RES1_O0;  //EXTERNAL
	output Tile_X11Y4_RES1_O1;  //EXTERNAL
	output Tile_X11Y4_RES1_O2;  //EXTERNAL
	output Tile_X11Y4_RES1_O3;  //EXTERNAL
	output Tile_X11Y4_RES2_O0;  //EXTERNAL
	output Tile_X11Y4_RES2_O1;  //EXTERNAL
	output Tile_X11Y4_RES2_O2;  //EXTERNAL
	output Tile_X11Y4_RES2_O3;  //EXTERNAL
	input Tile_X4Y5_OPA_I0;  //EXTERNAL
	input Tile_X4Y5_OPA_I1;  //EXTERNAL
	input Tile_X4Y5_OPA_I2;  //EXTERNAL
	input Tile_X4Y5_OPA_I3;  //EXTERNAL
	input Tile_X4Y5_OPB_I0;  //EXTERNAL
	input Tile_X4Y5_OPB_I1;  //EXTERNAL
	input Tile_X4Y5_OPB_I2;  //EXTERNAL
	input Tile_X4Y5_OPB_I3;  //EXTERNAL
	output Tile_X4Y5_RES0_O0;  //EXTERNAL
	output Tile_X4Y5_RES0_O1;  //EXTERNAL
	output Tile_X4Y5_RES0_O2;  //EXTERNAL
	output Tile_X4Y5_RES0_O3;  //EXTERNAL
	output Tile_X4Y5_RES1_O0;  //EXTERNAL
	output Tile_X4Y5_RES1_O1;  //EXTERNAL
	output Tile_X4Y5_RES1_O2;  //EXTERNAL
	output Tile_X4Y5_RES1_O3;  //EXTERNAL
	output Tile_X4Y5_RES2_O0;  //EXTERNAL
	output Tile_X4Y5_RES2_O1;  //EXTERNAL
	output Tile_X4Y5_RES2_O2;  //EXTERNAL
	output Tile_X4Y5_RES2_O3;  //EXTERNAL
	input Tile_X11Y5_OPA_I0;  //EXTERNAL
	input Tile_X11Y5_OPA_I1;  //EXTERNAL
	input Tile_X11Y5_OPA_I2;  //EXTERNAL
	input Tile_X11Y5_OPA_I3;  //EXTERNAL
	input Tile_X11Y5_OPB_I0;  //EXTERNAL
	input Tile_X11Y5_OPB_I1;  //EXTERNAL
	input Tile_X11Y5_OPB_I2;  //EXTERNAL
	input Tile_X11Y5_OPB_I3;  //EXTERNAL
	output Tile_X11Y5_RES0_O0;  //EXTERNAL
	output Tile_X11Y5_RES0_O1;  //EXTERNAL
	output Tile_X11Y5_RES0_O2;  //EXTERNAL
	output Tile_X11Y5_RES0_O3;  //EXTERNAL
	output Tile_X11Y5_RES1_O0;  //EXTERNAL
	output Tile_X11Y5_RES1_O1;  //EXTERNAL
	output Tile_X11Y5_RES1_O2;  //EXTERNAL
	output Tile_X11Y5_RES1_O3;  //EXTERNAL
	output Tile_X11Y5_RES2_O0;  //EXTERNAL
	output Tile_X11Y5_RES2_O1;  //EXTERNAL
	output Tile_X11Y5_RES2_O2;  //EXTERNAL
	output Tile_X11Y5_RES2_O3;  //EXTERNAL
	input Tile_X4Y6_OPA_I0;  //EXTERNAL
	input Tile_X4Y6_OPA_I1;  //EXTERNAL
	input Tile_X4Y6_OPA_I2;  //EXTERNAL
	input Tile_X4Y6_OPA_I3;  //EXTERNAL
	input Tile_X4Y6_OPB_I0;  //EXTERNAL
	input Tile_X4Y6_OPB_I1;  //EXTERNAL
	input Tile_X4Y6_OPB_I2;  //EXTERNAL
	input Tile_X4Y6_OPB_I3;  //EXTERNAL
	output Tile_X4Y6_RES0_O0;  //EXTERNAL
	output Tile_X4Y6_RES0_O1;  //EXTERNAL
	output Tile_X4Y6_RES0_O2;  //EXTERNAL
	output Tile_X4Y6_RES0_O3;  //EXTERNAL
	output Tile_X4Y6_RES1_O0;  //EXTERNAL
	output Tile_X4Y6_RES1_O1;  //EXTERNAL
	output Tile_X4Y6_RES1_O2;  //EXTERNAL
	output Tile_X4Y6_RES1_O3;  //EXTERNAL
	output Tile_X4Y6_RES2_O0;  //EXTERNAL
	output Tile_X4Y6_RES2_O1;  //EXTERNAL
	output Tile_X4Y6_RES2_O2;  //EXTERNAL
	output Tile_X4Y6_RES2_O3;  //EXTERNAL
	input Tile_X11Y6_OPA_I0;  //EXTERNAL
	input Tile_X11Y6_OPA_I1;  //EXTERNAL
	input Tile_X11Y6_OPA_I2;  //EXTERNAL
	input Tile_X11Y6_OPA_I3;  //EXTERNAL
	input Tile_X11Y6_OPB_I0;  //EXTERNAL
	input Tile_X11Y6_OPB_I1;  //EXTERNAL
	input Tile_X11Y6_OPB_I2;  //EXTERNAL
	input Tile_X11Y6_OPB_I3;  //EXTERNAL
	output Tile_X11Y6_RES0_O0;  //EXTERNAL
	output Tile_X11Y6_RES0_O1;  //EXTERNAL
	output Tile_X11Y6_RES0_O2;  //EXTERNAL
	output Tile_X11Y6_RES0_O3;  //EXTERNAL
	output Tile_X11Y6_RES1_O0;  //EXTERNAL
	output Tile_X11Y6_RES1_O1;  //EXTERNAL
	output Tile_X11Y6_RES1_O2;  //EXTERNAL
	output Tile_X11Y6_RES1_O3;  //EXTERNAL
	output Tile_X11Y6_RES2_O0;  //EXTERNAL
	output Tile_X11Y6_RES2_O1;  //EXTERNAL
	output Tile_X11Y6_RES2_O2;  //EXTERNAL
	output Tile_X11Y6_RES2_O3;  //EXTERNAL
	input Tile_X4Y7_OPA_I0;  //EXTERNAL
	input Tile_X4Y7_OPA_I1;  //EXTERNAL
	input Tile_X4Y7_OPA_I2;  //EXTERNAL
	input Tile_X4Y7_OPA_I3;  //EXTERNAL
	input Tile_X4Y7_OPB_I0;  //EXTERNAL
	input Tile_X4Y7_OPB_I1;  //EXTERNAL
	input Tile_X4Y7_OPB_I2;  //EXTERNAL
	input Tile_X4Y7_OPB_I3;  //EXTERNAL
	output Tile_X4Y7_RES0_O0;  //EXTERNAL
	output Tile_X4Y7_RES0_O1;  //EXTERNAL
	output Tile_X4Y7_RES0_O2;  //EXTERNAL
	output Tile_X4Y7_RES0_O3;  //EXTERNAL
	output Tile_X4Y7_RES1_O0;  //EXTERNAL
	output Tile_X4Y7_RES1_O1;  //EXTERNAL
	output Tile_X4Y7_RES1_O2;  //EXTERNAL
	output Tile_X4Y7_RES1_O3;  //EXTERNAL
	output Tile_X4Y7_RES2_O0;  //EXTERNAL
	output Tile_X4Y7_RES2_O1;  //EXTERNAL
	output Tile_X4Y7_RES2_O2;  //EXTERNAL
	output Tile_X4Y7_RES2_O3;  //EXTERNAL
	input Tile_X11Y7_OPA_I0;  //EXTERNAL
	input Tile_X11Y7_OPA_I1;  //EXTERNAL
	input Tile_X11Y7_OPA_I2;  //EXTERNAL
	input Tile_X11Y7_OPA_I3;  //EXTERNAL
	input Tile_X11Y7_OPB_I0;  //EXTERNAL
	input Tile_X11Y7_OPB_I1;  //EXTERNAL
	input Tile_X11Y7_OPB_I2;  //EXTERNAL
	input Tile_X11Y7_OPB_I3;  //EXTERNAL
	output Tile_X11Y7_RES0_O0;  //EXTERNAL
	output Tile_X11Y7_RES0_O1;  //EXTERNAL
	output Tile_X11Y7_RES0_O2;  //EXTERNAL
	output Tile_X11Y7_RES0_O3;  //EXTERNAL
	output Tile_X11Y7_RES1_O0;  //EXTERNAL
	output Tile_X11Y7_RES1_O1;  //EXTERNAL
	output Tile_X11Y7_RES1_O2;  //EXTERNAL
	output Tile_X11Y7_RES1_O3;  //EXTERNAL
	output Tile_X11Y7_RES2_O0;  //EXTERNAL
	output Tile_X11Y7_RES2_O1;  //EXTERNAL
	output Tile_X11Y7_RES2_O2;  //EXTERNAL
	output Tile_X11Y7_RES2_O3;  //EXTERNAL
	input Tile_X4Y8_OPA_I0;  //EXTERNAL
	input Tile_X4Y8_OPA_I1;  //EXTERNAL
	input Tile_X4Y8_OPA_I2;  //EXTERNAL
	input Tile_X4Y8_OPA_I3;  //EXTERNAL
	input Tile_X4Y8_OPB_I0;  //EXTERNAL
	input Tile_X4Y8_OPB_I1;  //EXTERNAL
	input Tile_X4Y8_OPB_I2;  //EXTERNAL
	input Tile_X4Y8_OPB_I3;  //EXTERNAL
	output Tile_X4Y8_RES0_O0;  //EXTERNAL
	output Tile_X4Y8_RES0_O1;  //EXTERNAL
	output Tile_X4Y8_RES0_O2;  //EXTERNAL
	output Tile_X4Y8_RES0_O3;  //EXTERNAL
	output Tile_X4Y8_RES1_O0;  //EXTERNAL
	output Tile_X4Y8_RES1_O1;  //EXTERNAL
	output Tile_X4Y8_RES1_O2;  //EXTERNAL
	output Tile_X4Y8_RES1_O3;  //EXTERNAL
	output Tile_X4Y8_RES2_O0;  //EXTERNAL
	output Tile_X4Y8_RES2_O1;  //EXTERNAL
	output Tile_X4Y8_RES2_O2;  //EXTERNAL
	output Tile_X4Y8_RES2_O3;  //EXTERNAL
	input Tile_X11Y8_OPA_I0;  //EXTERNAL
	input Tile_X11Y8_OPA_I1;  //EXTERNAL
	input Tile_X11Y8_OPA_I2;  //EXTERNAL
	input Tile_X11Y8_OPA_I3;  //EXTERNAL
	input Tile_X11Y8_OPB_I0;  //EXTERNAL
	input Tile_X11Y8_OPB_I1;  //EXTERNAL
	input Tile_X11Y8_OPB_I2;  //EXTERNAL
	input Tile_X11Y8_OPB_I3;  //EXTERNAL
	output Tile_X11Y8_RES0_O0;  //EXTERNAL
	output Tile_X11Y8_RES0_O1;  //EXTERNAL
	output Tile_X11Y8_RES0_O2;  //EXTERNAL
	output Tile_X11Y8_RES0_O3;  //EXTERNAL
	output Tile_X11Y8_RES1_O0;  //EXTERNAL
	output Tile_X11Y8_RES1_O1;  //EXTERNAL
	output Tile_X11Y8_RES1_O2;  //EXTERNAL
	output Tile_X11Y8_RES1_O3;  //EXTERNAL
	output Tile_X11Y8_RES2_O0;  //EXTERNAL
	output Tile_X11Y8_RES2_O1;  //EXTERNAL
	output Tile_X11Y8_RES2_O2;  //EXTERNAL
	output Tile_X11Y8_RES2_O3;  //EXTERNAL
	input Tile_X4Y9_OPA_I0;  //EXTERNAL
	input Tile_X4Y9_OPA_I1;  //EXTERNAL
	input Tile_X4Y9_OPA_I2;  //EXTERNAL
	input Tile_X4Y9_OPA_I3;  //EXTERNAL
	input Tile_X4Y9_OPB_I0;  //EXTERNAL
	input Tile_X4Y9_OPB_I1;  //EXTERNAL
	input Tile_X4Y9_OPB_I2;  //EXTERNAL
	input Tile_X4Y9_OPB_I3;  //EXTERNAL
	output Tile_X4Y9_RES0_O0;  //EXTERNAL
	output Tile_X4Y9_RES0_O1;  //EXTERNAL
	output Tile_X4Y9_RES0_O2;  //EXTERNAL
	output Tile_X4Y9_RES0_O3;  //EXTERNAL
	output Tile_X4Y9_RES1_O0;  //EXTERNAL
	output Tile_X4Y9_RES1_O1;  //EXTERNAL
	output Tile_X4Y9_RES1_O2;  //EXTERNAL
	output Tile_X4Y9_RES1_O3;  //EXTERNAL
	output Tile_X4Y9_RES2_O0;  //EXTERNAL
	output Tile_X4Y9_RES2_O1;  //EXTERNAL
	output Tile_X4Y9_RES2_O2;  //EXTERNAL
	output Tile_X4Y9_RES2_O3;  //EXTERNAL
	input Tile_X11Y9_OPA_I0;  //EXTERNAL
	input Tile_X11Y9_OPA_I1;  //EXTERNAL
	input Tile_X11Y9_OPA_I2;  //EXTERNAL
	input Tile_X11Y9_OPA_I3;  //EXTERNAL
	input Tile_X11Y9_OPB_I0;  //EXTERNAL
	input Tile_X11Y9_OPB_I1;  //EXTERNAL
	input Tile_X11Y9_OPB_I2;  //EXTERNAL
	input Tile_X11Y9_OPB_I3;  //EXTERNAL
	output Tile_X11Y9_RES0_O0;  //EXTERNAL
	output Tile_X11Y9_RES0_O1;  //EXTERNAL
	output Tile_X11Y9_RES0_O2;  //EXTERNAL
	output Tile_X11Y9_RES0_O3;  //EXTERNAL
	output Tile_X11Y9_RES1_O0;  //EXTERNAL
	output Tile_X11Y9_RES1_O1;  //EXTERNAL
	output Tile_X11Y9_RES1_O2;  //EXTERNAL
	output Tile_X11Y9_RES1_O3;  //EXTERNAL
	output Tile_X11Y9_RES2_O0;  //EXTERNAL
	output Tile_X11Y9_RES2_O1;  //EXTERNAL
	output Tile_X11Y9_RES2_O2;  //EXTERNAL
	output Tile_X11Y9_RES2_O3;  //EXTERNAL
	output Tile_X0Y10_A_I_top;   //EXTERNAL has to ge to top-level entity not the switch matrix
	output Tile_X0Y10_A_T_top;   //EXTERNAL has to ge to top-level entity not the switch matrix
	input Tile_X0Y10_A_O_top;   //EXTERNAL has to ge to top-level entity not the switch matrix
	output Tile_X0Y10_B_I_top;   //EXTERNAL has to ge to top-level entity not the switch matrix
	output Tile_X0Y10_B_T_top;   //EXTERNAL has to ge to top-level entity not the switch matrix
	input Tile_X0Y10_B_O_top;   //EXTERNAL has to ge to top-level entity not the switch matrix
	output Tile_X0Y10_A_config_C_bit0;  //EXTERNAL
	output Tile_X0Y10_A_config_C_bit1;  //EXTERNAL
	output Tile_X0Y10_A_config_C_bit2;  //EXTERNAL
	output Tile_X0Y10_A_config_C_bit3;  //EXTERNAL
	output Tile_X0Y10_B_config_C_bit0;  //EXTERNAL
	output Tile_X0Y10_B_config_C_bit1;  //EXTERNAL
	output Tile_X0Y10_B_config_C_bit2;  //EXTERNAL
	output Tile_X0Y10_B_config_C_bit3;  //EXTERNAL
	input Tile_X15Y10_RAM2FAB_D0_I0;  //EXTERNAL
	input Tile_X15Y10_RAM2FAB_D0_I1;  //EXTERNAL
	input Tile_X15Y10_RAM2FAB_D0_I2;  //EXTERNAL
	input Tile_X15Y10_RAM2FAB_D0_I3;  //EXTERNAL
	input Tile_X15Y10_RAM2FAB_D1_I0;  //EXTERNAL
	input Tile_X15Y10_RAM2FAB_D1_I1;  //EXTERNAL
	input Tile_X15Y10_RAM2FAB_D1_I2;  //EXTERNAL
	input Tile_X15Y10_RAM2FAB_D1_I3;  //EXTERNAL
	input Tile_X15Y10_RAM2FAB_D2_I0;  //EXTERNAL
	input Tile_X15Y10_RAM2FAB_D2_I1;  //EXTERNAL
	input Tile_X15Y10_RAM2FAB_D2_I2;  //EXTERNAL
	input Tile_X15Y10_RAM2FAB_D2_I3;  //EXTERNAL
	input Tile_X15Y10_RAM2FAB_D3_I0;  //EXTERNAL
	input Tile_X15Y10_RAM2FAB_D3_I1;  //EXTERNAL
	input Tile_X15Y10_RAM2FAB_D3_I2;  //EXTERNAL
	input Tile_X15Y10_RAM2FAB_D3_I3;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_D0_O0;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_D0_O1;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_D0_O2;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_D0_O3;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_D1_O0;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_D1_O1;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_D1_O2;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_D1_O3;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_D2_O0;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_D2_O1;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_D2_O2;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_D2_O3;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_D3_O0;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_D3_O1;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_D3_O2;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_D3_O3;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_A0_O0;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_A0_O1;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_A0_O2;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_A0_O3;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_A1_O0;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_A1_O1;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_A1_O2;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_A1_O3;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_C_O0;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_C_O1;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_C_O2;  //EXTERNAL
	output Tile_X15Y10_FAB2RAM_C_O3;  //EXTERNAL
	output Tile_X15Y10_Config_accessC_bit0;  //EXTERNAL
	output Tile_X15Y10_Config_accessC_bit1;  //EXTERNAL
	output Tile_X15Y10_Config_accessC_bit2;  //EXTERNAL
	output Tile_X15Y10_Config_accessC_bit3;  //EXTERNAL
	output Tile_X0Y11_A_I_top;   //EXTERNAL has to ge to top-level entity not the switch matrix
	output Tile_X0Y11_A_T_top;   //EXTERNAL has to ge to top-level entity not the switch matrix
	input Tile_X0Y11_A_O_top;   //EXTERNAL has to ge to top-level entity not the switch matrix
	output Tile_X0Y11_B_I_top;   //EXTERNAL has to ge to top-level entity not the switch matrix
	output Tile_X0Y11_B_T_top;   //EXTERNAL has to ge to top-level entity not the switch matrix
	input Tile_X0Y11_B_O_top;   //EXTERNAL has to ge to top-level entity not the switch matrix
	output Tile_X0Y11_A_config_C_bit0;  //EXTERNAL
	output Tile_X0Y11_A_config_C_bit1;  //EXTERNAL
	output Tile_X0Y11_A_config_C_bit2;  //EXTERNAL
	output Tile_X0Y11_A_config_C_bit3;  //EXTERNAL
	output Tile_X0Y11_B_config_C_bit0;  //EXTERNAL
	output Tile_X0Y11_B_config_C_bit1;  //EXTERNAL
	output Tile_X0Y11_B_config_C_bit2;  //EXTERNAL
	output Tile_X0Y11_B_config_C_bit3;  //EXTERNAL
	input Tile_X15Y11_RAM2FAB_D0_I0;  //EXTERNAL
	input Tile_X15Y11_RAM2FAB_D0_I1;  //EXTERNAL
	input Tile_X15Y11_RAM2FAB_D0_I2;  //EXTERNAL
	input Tile_X15Y11_RAM2FAB_D0_I3;  //EXTERNAL
	input Tile_X15Y11_RAM2FAB_D1_I0;  //EXTERNAL
	input Tile_X15Y11_RAM2FAB_D1_I1;  //EXTERNAL
	input Tile_X15Y11_RAM2FAB_D1_I2;  //EXTERNAL
	input Tile_X15Y11_RAM2FAB_D1_I3;  //EXTERNAL
	input Tile_X15Y11_RAM2FAB_D2_I0;  //EXTERNAL
	input Tile_X15Y11_RAM2FAB_D2_I1;  //EXTERNAL
	input Tile_X15Y11_RAM2FAB_D2_I2;  //EXTERNAL
	input Tile_X15Y11_RAM2FAB_D2_I3;  //EXTERNAL
	input Tile_X15Y11_RAM2FAB_D3_I0;  //EXTERNAL
	input Tile_X15Y11_RAM2FAB_D3_I1;  //EXTERNAL
	input Tile_X15Y11_RAM2FAB_D3_I2;  //EXTERNAL
	input Tile_X15Y11_RAM2FAB_D3_I3;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_D0_O0;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_D0_O1;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_D0_O2;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_D0_O3;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_D1_O0;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_D1_O1;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_D1_O2;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_D1_O3;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_D2_O0;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_D2_O1;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_D2_O2;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_D2_O3;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_D3_O0;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_D3_O1;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_D3_O2;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_D3_O3;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_A0_O0;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_A0_O1;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_A0_O2;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_A0_O3;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_A1_O0;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_A1_O1;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_A1_O2;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_A1_O3;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_C_O0;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_C_O1;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_C_O2;  //EXTERNAL
	output Tile_X15Y11_FAB2RAM_C_O3;  //EXTERNAL
	output Tile_X15Y11_Config_accessC_bit0;  //EXTERNAL
	output Tile_X15Y11_Config_accessC_bit1;  //EXTERNAL
	output Tile_X15Y11_Config_accessC_bit2;  //EXTERNAL
	output Tile_X15Y11_Config_accessC_bit3;  //EXTERNAL
	output Tile_X0Y12_A_I_top;   //EXTERNAL has to ge to top-level entity not the switch matrix
	output Tile_X0Y12_A_T_top;   //EXTERNAL has to ge to top-level entity not the switch matrix
	input Tile_X0Y12_A_O_top;   //EXTERNAL has to ge to top-level entity not the switch matrix
	output Tile_X0Y12_B_I_top;   //EXTERNAL has to ge to top-level entity not the switch matrix
	output Tile_X0Y12_B_T_top;   //EXTERNAL has to ge to top-level entity not the switch matrix
	input Tile_X0Y12_B_O_top;   //EXTERNAL has to ge to top-level entity not the switch matrix
	output Tile_X0Y12_A_config_C_bit0;  //EXTERNAL
	output Tile_X0Y12_A_config_C_bit1;  //EXTERNAL
	output Tile_X0Y12_A_config_C_bit2;  //EXTERNAL
	output Tile_X0Y12_A_config_C_bit3;  //EXTERNAL
	output Tile_X0Y12_B_config_C_bit0;  //EXTERNAL
	output Tile_X0Y12_B_config_C_bit1;  //EXTERNAL
	output Tile_X0Y12_B_config_C_bit2;  //EXTERNAL
	output Tile_X0Y12_B_config_C_bit3;  //EXTERNAL
	input Tile_X15Y12_RAM2FAB_D0_I0;  //EXTERNAL
	input Tile_X15Y12_RAM2FAB_D0_I1;  //EXTERNAL
	input Tile_X15Y12_RAM2FAB_D0_I2;  //EXTERNAL
	input Tile_X15Y12_RAM2FAB_D0_I3;  //EXTERNAL
	input Tile_X15Y12_RAM2FAB_D1_I0;  //EXTERNAL
	input Tile_X15Y12_RAM2FAB_D1_I1;  //EXTERNAL
	input Tile_X15Y12_RAM2FAB_D1_I2;  //EXTERNAL
	input Tile_X15Y12_RAM2FAB_D1_I3;  //EXTERNAL
	input Tile_X15Y12_RAM2FAB_D2_I0;  //EXTERNAL
	input Tile_X15Y12_RAM2FAB_D2_I1;  //EXTERNAL
	input Tile_X15Y12_RAM2FAB_D2_I2;  //EXTERNAL
	input Tile_X15Y12_RAM2FAB_D2_I3;  //EXTERNAL
	input Tile_X15Y12_RAM2FAB_D3_I0;  //EXTERNAL
	input Tile_X15Y12_RAM2FAB_D3_I1;  //EXTERNAL
	input Tile_X15Y12_RAM2FAB_D3_I2;  //EXTERNAL
	input Tile_X15Y12_RAM2FAB_D3_I3;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_D0_O0;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_D0_O1;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_D0_O2;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_D0_O3;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_D1_O0;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_D1_O1;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_D1_O2;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_D1_O3;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_D2_O0;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_D2_O1;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_D2_O2;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_D2_O3;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_D3_O0;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_D3_O1;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_D3_O2;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_D3_O3;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_A0_O0;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_A0_O1;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_A0_O2;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_A0_O3;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_A1_O0;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_A1_O1;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_A1_O2;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_A1_O3;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_C_O0;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_C_O1;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_C_O2;  //EXTERNAL
	output Tile_X15Y12_FAB2RAM_C_O3;  //EXTERNAL
	output Tile_X15Y12_Config_accessC_bit0;  //EXTERNAL
	output Tile_X15Y12_Config_accessC_bit1;  //EXTERNAL
	output Tile_X15Y12_Config_accessC_bit2;  //EXTERNAL
	output Tile_X15Y12_Config_accessC_bit3;  //EXTERNAL
	input [(FrameBitsPerRow*14)-1:0] FrameData;   // CONFIG_PORT this is a keyword needed to connect the tile to the bitstream frame register
	input [(MaxFramesPerCol*16)-1:0] FrameStrobe;   // CONFIG_PORT this is a keyword needed to connect the tile to the bitstream frame register 
	//global


//signal declarations
	wire Tile_X0Y0_UserCLKo;
	wire Tile_X1Y0_UserCLKo;
	wire Tile_X2Y0_UserCLKo;
	wire Tile_X3Y0_UserCLKo;
	wire Tile_X4Y0_UserCLKo;
	wire Tile_X5Y0_UserCLKo;
	wire Tile_X6Y0_UserCLKo;
	wire Tile_X7Y0_UserCLKo;
	wire Tile_X8Y0_UserCLKo;
	wire Tile_X9Y0_UserCLKo;
	wire Tile_X10Y0_UserCLKo;
	wire Tile_X11Y0_UserCLKo;
	wire Tile_X12Y0_UserCLKo;
	wire Tile_X13Y0_UserCLKo;
	wire Tile_X14Y0_UserCLKo;
	wire Tile_X15Y0_UserCLKo;
	wire Tile_X0Y1_UserCLKo;
	wire Tile_X1Y1_UserCLKo;
	wire Tile_X2Y1_UserCLKo;
	wire Tile_X3Y1_UserCLKo;
	wire Tile_X4Y1_UserCLKo;
	wire Tile_X5Y1_UserCLKo;
	wire Tile_X6Y1_UserCLKo;
	wire Tile_X7Y1_UserCLKo;
	wire Tile_X8Y1_UserCLKo;
	wire Tile_X9Y1_UserCLKo;
	wire Tile_X10Y1_UserCLKo;
	wire Tile_X11Y1_UserCLKo;
	wire Tile_X12Y1_UserCLKo;
	wire Tile_X13Y1_UserCLKo;
	wire Tile_X14Y1_UserCLKo;
	wire Tile_X15Y1_UserCLKo;
	wire Tile_X0Y2_UserCLKo;
	wire Tile_X1Y2_UserCLKo;
	wire Tile_X2Y2_UserCLKo;
	wire Tile_X3Y2_UserCLKo;
	wire Tile_X4Y2_UserCLKo;
	wire Tile_X5Y2_UserCLKo;
	wire Tile_X6Y2_UserCLKo;
	wire Tile_X7Y2_UserCLKo;
	wire Tile_X8Y2_UserCLKo;
	wire Tile_X9Y2_UserCLKo;
	wire Tile_X10Y2_UserCLKo;
	wire Tile_X11Y2_UserCLKo;
	wire Tile_X12Y2_UserCLKo;
	wire Tile_X13Y2_UserCLKo;
	wire Tile_X14Y2_UserCLKo;
	wire Tile_X15Y2_UserCLKo;
	wire Tile_X0Y3_UserCLKo;
	wire Tile_X1Y3_UserCLKo;
	wire Tile_X2Y3_UserCLKo;
	wire Tile_X3Y3_UserCLKo;
	wire Tile_X4Y3_UserCLKo;
	wire Tile_X5Y3_UserCLKo;
	wire Tile_X6Y3_UserCLKo;
	wire Tile_X7Y3_UserCLKo;
	wire Tile_X8Y3_UserCLKo;
	wire Tile_X9Y3_UserCLKo;
	wire Tile_X10Y3_UserCLKo;
	wire Tile_X11Y3_UserCLKo;
	wire Tile_X12Y3_UserCLKo;
	wire Tile_X13Y3_UserCLKo;
	wire Tile_X14Y3_UserCLKo;
	wire Tile_X15Y3_UserCLKo;
	wire Tile_X0Y4_UserCLKo;
	wire Tile_X1Y4_UserCLKo;
	wire Tile_X2Y4_UserCLKo;
	wire Tile_X3Y4_UserCLKo;
	wire Tile_X4Y4_UserCLKo;
	wire Tile_X5Y4_UserCLKo;
	wire Tile_X6Y4_UserCLKo;
	wire Tile_X7Y4_UserCLKo;
	wire Tile_X8Y4_UserCLKo;
	wire Tile_X9Y4_UserCLKo;
	wire Tile_X10Y4_UserCLKo;
	wire Tile_X11Y4_UserCLKo;
	wire Tile_X12Y4_UserCLKo;
	wire Tile_X13Y4_UserCLKo;
	wire Tile_X14Y4_UserCLKo;
	wire Tile_X15Y4_UserCLKo;
	wire Tile_X0Y5_UserCLKo;
	wire Tile_X1Y5_UserCLKo;
	wire Tile_X2Y5_UserCLKo;
	wire Tile_X3Y5_UserCLKo;
	wire Tile_X4Y5_UserCLKo;
	wire Tile_X5Y5_UserCLKo;
	wire Tile_X6Y5_UserCLKo;
	wire Tile_X7Y5_UserCLKo;
	wire Tile_X8Y5_UserCLKo;
	wire Tile_X9Y5_UserCLKo;
	wire Tile_X10Y5_UserCLKo;
	wire Tile_X11Y5_UserCLKo;
	wire Tile_X12Y5_UserCLKo;
	wire Tile_X13Y5_UserCLKo;
	wire Tile_X14Y5_UserCLKo;
	wire Tile_X15Y5_UserCLKo;
	wire Tile_X0Y6_UserCLKo;
	wire Tile_X1Y6_UserCLKo;
	wire Tile_X2Y6_UserCLKo;
	wire Tile_X3Y6_UserCLKo;
	wire Tile_X4Y6_UserCLKo;
	wire Tile_X5Y6_UserCLKo;
	wire Tile_X6Y6_UserCLKo;
	wire Tile_X7Y6_UserCLKo;
	wire Tile_X8Y6_UserCLKo;
	wire Tile_X9Y6_UserCLKo;
	wire Tile_X10Y6_UserCLKo;
	wire Tile_X11Y6_UserCLKo;
	wire Tile_X12Y6_UserCLKo;
	wire Tile_X13Y6_UserCLKo;
	wire Tile_X14Y6_UserCLKo;
	wire Tile_X15Y6_UserCLKo;
	wire Tile_X0Y7_UserCLKo;
	wire Tile_X1Y7_UserCLKo;
	wire Tile_X2Y7_UserCLKo;
	wire Tile_X3Y7_UserCLKo;
	wire Tile_X4Y7_UserCLKo;
	wire Tile_X5Y7_UserCLKo;
	wire Tile_X6Y7_UserCLKo;
	wire Tile_X7Y7_UserCLKo;
	wire Tile_X8Y7_UserCLKo;
	wire Tile_X9Y7_UserCLKo;
	wire Tile_X10Y7_UserCLKo;
	wire Tile_X11Y7_UserCLKo;
	wire Tile_X12Y7_UserCLKo;
	wire Tile_X13Y7_UserCLKo;
	wire Tile_X14Y7_UserCLKo;
	wire Tile_X15Y7_UserCLKo;
	wire Tile_X0Y8_UserCLKo;
	wire Tile_X1Y8_UserCLKo;
	wire Tile_X2Y8_UserCLKo;
	wire Tile_X3Y8_UserCLKo;
	wire Tile_X4Y8_UserCLKo;
	wire Tile_X5Y8_UserCLKo;
	wire Tile_X6Y8_UserCLKo;
	wire Tile_X7Y8_UserCLKo;
	wire Tile_X8Y8_UserCLKo;
	wire Tile_X9Y8_UserCLKo;
	wire Tile_X10Y8_UserCLKo;
	wire Tile_X11Y8_UserCLKo;
	wire Tile_X12Y8_UserCLKo;
	wire Tile_X13Y8_UserCLKo;
	wire Tile_X14Y8_UserCLKo;
	wire Tile_X15Y8_UserCLKo;
	wire Tile_X0Y9_UserCLKo;
	wire Tile_X1Y9_UserCLKo;
	wire Tile_X2Y9_UserCLKo;
	wire Tile_X3Y9_UserCLKo;
	wire Tile_X4Y9_UserCLKo;
	wire Tile_X5Y9_UserCLKo;
	wire Tile_X6Y9_UserCLKo;
	wire Tile_X7Y9_UserCLKo;
	wire Tile_X8Y9_UserCLKo;
	wire Tile_X9Y9_UserCLKo;
	wire Tile_X10Y9_UserCLKo;
	wire Tile_X11Y9_UserCLKo;
	wire Tile_X12Y9_UserCLKo;
	wire Tile_X13Y9_UserCLKo;
	wire Tile_X14Y9_UserCLKo;
	wire Tile_X15Y9_UserCLKo;
	wire Tile_X0Y10_UserCLKo;
	wire Tile_X1Y10_UserCLKo;
	wire Tile_X2Y10_UserCLKo;
	wire Tile_X3Y10_UserCLKo;
	wire Tile_X4Y10_UserCLKo;
	wire Tile_X5Y10_UserCLKo;
	wire Tile_X6Y10_UserCLKo;
	wire Tile_X7Y10_UserCLKo;
	wire Tile_X8Y10_UserCLKo;
	wire Tile_X9Y10_UserCLKo;
	wire Tile_X10Y10_UserCLKo;
	wire Tile_X11Y10_UserCLKo;
	wire Tile_X12Y10_UserCLKo;
	wire Tile_X13Y10_UserCLKo;
	wire Tile_X14Y10_UserCLKo;
	wire Tile_X15Y10_UserCLKo;
	wire Tile_X0Y11_UserCLKo;
	wire Tile_X1Y11_UserCLKo;
	wire Tile_X2Y11_UserCLKo;
	wire Tile_X3Y11_UserCLKo;
	wire Tile_X4Y11_UserCLKo;
	wire Tile_X5Y11_UserCLKo;
	wire Tile_X6Y11_UserCLKo;
	wire Tile_X7Y11_UserCLKo;
	wire Tile_X8Y11_UserCLKo;
	wire Tile_X9Y11_UserCLKo;
	wire Tile_X10Y11_UserCLKo;
	wire Tile_X11Y11_UserCLKo;
	wire Tile_X12Y11_UserCLKo;
	wire Tile_X13Y11_UserCLKo;
	wire Tile_X14Y11_UserCLKo;
	wire Tile_X15Y11_UserCLKo;
	wire Tile_X0Y12_UserCLKo;
	wire Tile_X1Y12_UserCLKo;
	wire Tile_X2Y12_UserCLKo;
	wire Tile_X3Y12_UserCLKo;
	wire Tile_X4Y12_UserCLKo;
	wire Tile_X5Y12_UserCLKo;
	wire Tile_X6Y12_UserCLKo;
	wire Tile_X7Y12_UserCLKo;
	wire Tile_X8Y12_UserCLKo;
	wire Tile_X9Y12_UserCLKo;
	wire Tile_X10Y12_UserCLKo;
	wire Tile_X11Y12_UserCLKo;
	wire Tile_X12Y12_UserCLKo;
	wire Tile_X13Y12_UserCLKo;
	wire Tile_X14Y12_UserCLKo;
	wire Tile_X15Y12_UserCLKo;
	wire Tile_X0Y13_UserCLKo;
	wire Tile_X1Y13_UserCLKo;
	wire Tile_X2Y13_UserCLKo;
	wire Tile_X3Y13_UserCLKo;
	wire Tile_X4Y13_UserCLKo;
	wire Tile_X5Y13_UserCLKo;
	wire Tile_X6Y13_UserCLKo;
	wire Tile_X7Y13_UserCLKo;
	wire Tile_X8Y13_UserCLKo;
	wire Tile_X9Y13_UserCLKo;
	wire Tile_X10Y13_UserCLKo;
	wire Tile_X11Y13_UserCLKo;
	wire Tile_X12Y13_UserCLKo;
	wire Tile_X13Y13_UserCLKo;
	wire Tile_X14Y13_UserCLKo;
	wire Tile_X15Y13_UserCLKo;
//configuration signal declarations

	wire [FrameBitsPerRow-1:0] Tile_Y1_FrameData;
	wire [FrameBitsPerRow-1:0] Tile_Y2_FrameData;
	wire [FrameBitsPerRow-1:0] Tile_Y3_FrameData;
	wire [FrameBitsPerRow-1:0] Tile_Y4_FrameData;
	wire [FrameBitsPerRow-1:0] Tile_Y5_FrameData;
	wire [FrameBitsPerRow-1:0] Tile_Y6_FrameData;
	wire [FrameBitsPerRow-1:0] Tile_Y7_FrameData;
	wire [FrameBitsPerRow-1:0] Tile_Y8_FrameData;
	wire [FrameBitsPerRow-1:0] Tile_Y9_FrameData;
	wire [FrameBitsPerRow-1:0] Tile_Y10_FrameData;
	wire [FrameBitsPerRow-1:0] Tile_Y11_FrameData;
	wire [FrameBitsPerRow-1:0] Tile_Y12_FrameData;
	wire [MaxFramesPerCol-1:0] Tile_X0_FrameStrobe;
	wire [MaxFramesPerCol-1:0] Tile_X1_FrameStrobe;
	wire [MaxFramesPerCol-1:0] Tile_X2_FrameStrobe;
	wire [MaxFramesPerCol-1:0] Tile_X3_FrameStrobe;
	wire [MaxFramesPerCol-1:0] Tile_X4_FrameStrobe;
	wire [MaxFramesPerCol-1:0] Tile_X5_FrameStrobe;
	wire [MaxFramesPerCol-1:0] Tile_X6_FrameStrobe;
	wire [MaxFramesPerCol-1:0] Tile_X7_FrameStrobe;
	wire [MaxFramesPerCol-1:0] Tile_X8_FrameStrobe;
	wire [MaxFramesPerCol-1:0] Tile_X9_FrameStrobe;
	wire [MaxFramesPerCol-1:0] Tile_X10_FrameStrobe;
	wire [MaxFramesPerCol-1:0] Tile_X11_FrameStrobe;
	wire [MaxFramesPerCol-1:0] Tile_X12_FrameStrobe;
	wire [MaxFramesPerCol-1:0] Tile_X13_FrameStrobe;
	wire [MaxFramesPerCol-1:0] Tile_X14_FrameStrobe;
	wire [MaxFramesPerCol-1:0] Tile_X15_FrameStrobe;
	wire [FrameBitsPerRow-1:0] Tile_X0Y1_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X1Y1_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X2Y1_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X3Y1_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X4Y1_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X5Y1_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X6Y1_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X7Y1_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X8Y1_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X9Y1_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X10Y1_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X11Y1_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X12Y1_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X13Y1_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X14Y1_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X15Y1_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X0Y2_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X1Y2_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X2Y2_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X3Y2_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X4Y2_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X5Y2_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X6Y2_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X7Y2_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X8Y2_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X9Y2_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X10Y2_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X11Y2_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X12Y2_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X13Y2_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X14Y2_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X15Y2_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X0Y3_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X1Y3_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X2Y3_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X3Y3_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X4Y3_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X5Y3_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X6Y3_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X7Y3_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X8Y3_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X9Y3_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X10Y3_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X11Y3_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X12Y3_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X13Y3_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X14Y3_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X15Y3_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X0Y4_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X1Y4_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X2Y4_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X3Y4_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X4Y4_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X5Y4_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X6Y4_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X7Y4_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X8Y4_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X9Y4_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X10Y4_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X11Y4_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X12Y4_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X13Y4_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X14Y4_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X15Y4_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X0Y5_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X1Y5_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X2Y5_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X3Y5_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X4Y5_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X5Y5_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X6Y5_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X7Y5_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X8Y5_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X9Y5_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X10Y5_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X11Y5_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X12Y5_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X13Y5_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X14Y5_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X15Y5_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X0Y6_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X1Y6_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X2Y6_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X3Y6_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X4Y6_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X5Y6_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X6Y6_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X7Y6_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X8Y6_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X9Y6_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X10Y6_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X11Y6_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X12Y6_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X13Y6_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X14Y6_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X15Y6_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X0Y7_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X1Y7_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X2Y7_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X3Y7_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X4Y7_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X5Y7_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X6Y7_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X7Y7_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X8Y7_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X9Y7_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X10Y7_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X11Y7_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X12Y7_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X13Y7_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X14Y7_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X15Y7_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X0Y8_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X1Y8_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X2Y8_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X3Y8_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X4Y8_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X5Y8_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X6Y8_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X7Y8_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X8Y8_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X9Y8_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X10Y8_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X11Y8_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X12Y8_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X13Y8_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X14Y8_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X15Y8_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X0Y9_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X1Y9_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X2Y9_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X3Y9_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X4Y9_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X5Y9_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X6Y9_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X7Y9_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X8Y9_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X9Y9_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X10Y9_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X11Y9_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X12Y9_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X13Y9_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X14Y9_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X15Y9_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X0Y10_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X1Y10_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X2Y10_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X3Y10_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X4Y10_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X5Y10_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X6Y10_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X7Y10_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X8Y10_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X9Y10_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X10Y10_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X11Y10_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X12Y10_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X13Y10_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X14Y10_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X15Y10_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X0Y11_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X1Y11_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X2Y11_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X3Y11_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X4Y11_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X5Y11_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X6Y11_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X7Y11_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X8Y11_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X9Y11_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X10Y11_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X11Y11_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X12Y11_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X13Y11_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X14Y11_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X15Y11_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X0Y12_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X1Y12_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X2Y12_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X3Y12_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X4Y12_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X5Y12_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X6Y12_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X7Y12_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X8Y12_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X9Y12_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X10Y12_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X11Y12_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X12Y12_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X13Y12_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X14Y12_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X15Y12_FrameData_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y0_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y0_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y0_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y0_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y0_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y0_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y0_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y0_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X8Y0_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X9Y0_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X10Y0_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X11Y0_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X12Y0_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X13Y0_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X14Y0_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X15Y0_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y1_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y1_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y1_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y1_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y1_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y1_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y1_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y1_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X8Y1_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X9Y1_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X10Y1_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X11Y1_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X12Y1_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X13Y1_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X14Y1_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X15Y1_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y2_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y2_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y2_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y2_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y2_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y2_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y2_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y2_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X8Y2_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X9Y2_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X10Y2_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X11Y2_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X12Y2_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X13Y2_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X14Y2_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X15Y2_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y3_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y3_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y3_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y3_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y3_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y3_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y3_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y3_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X8Y3_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X9Y3_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X10Y3_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X11Y3_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X12Y3_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X13Y3_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X14Y3_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X15Y3_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y4_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y4_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y4_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y4_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y4_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y4_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y4_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y4_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X8Y4_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X9Y4_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X10Y4_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X11Y4_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X12Y4_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X13Y4_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X14Y4_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X15Y4_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y5_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y5_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y5_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y5_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y5_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y5_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y5_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y5_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X8Y5_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X9Y5_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X10Y5_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X11Y5_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X12Y5_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X13Y5_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X14Y5_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X15Y5_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y6_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y6_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y6_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y6_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y6_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y6_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y6_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y6_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X8Y6_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X9Y6_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X10Y6_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X11Y6_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X12Y6_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X13Y6_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X14Y6_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X15Y6_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y7_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y7_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y7_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y7_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y7_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y7_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y7_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y7_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X8Y7_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X9Y7_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X10Y7_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X11Y7_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X12Y7_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X13Y7_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X14Y7_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X15Y7_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y8_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y8_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y8_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y8_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y8_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y8_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y8_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y8_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X8Y8_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X9Y8_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X10Y8_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X11Y8_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X12Y8_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X13Y8_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X14Y8_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X15Y8_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y9_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y9_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y9_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y9_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y9_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y9_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y9_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y9_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X8Y9_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X9Y9_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X10Y9_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X11Y9_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X12Y9_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X13Y9_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X14Y9_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X15Y9_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y10_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y10_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y10_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y10_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y10_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y10_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y10_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y10_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X8Y10_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X9Y10_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X10Y10_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X11Y10_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X12Y10_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X13Y10_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X14Y10_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X15Y10_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y11_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y11_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y11_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y11_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y11_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y11_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y11_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y11_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X8Y11_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X9Y11_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X10Y11_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X11Y11_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X12Y11_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X13Y11_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X14Y11_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X15Y11_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y12_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y12_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y12_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y12_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y12_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y12_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y12_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y12_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X8Y12_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X9Y12_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X10Y12_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X11Y12_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X12Y12_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X13Y12_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X14Y12_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X15Y12_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y13_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y13_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y13_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y13_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y13_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y13_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y13_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y13_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X8Y13_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X9Y13_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X10Y13_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X11Y13_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X12Y13_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X13Y13_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X14Y13_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X15Y13_FrameStrobe_O;

//tile-to-tile signal declarations

	wire [3:0] Tile_X5Y0_S1BEG;
	wire [7:0] Tile_X5Y0_S2BEG;
	wire [7:0] Tile_X5Y0_S2BEGb;
	wire [15:0] Tile_X5Y0_S4BEG;
	wire [15:0] Tile_X5Y0_SS4BEG;
	wire [3:0] Tile_X6Y0_S1BEG;
	wire [7:0] Tile_X6Y0_S2BEG;
	wire [7:0] Tile_X6Y0_S2BEGb;
	wire [15:0] Tile_X6Y0_S4BEG;
	wire [15:0] Tile_X6Y0_SS4BEG;
	wire [3:0] Tile_X7Y0_S1BEG;
	wire [7:0] Tile_X7Y0_S2BEG;
	wire [7:0] Tile_X7Y0_S2BEGb;
	wire [15:0] Tile_X7Y0_S4BEG;
	wire [15:0] Tile_X7Y0_SS4BEG;
	wire [3:0] Tile_X8Y0_S1BEG;
	wire [7:0] Tile_X8Y0_S2BEG;
	wire [7:0] Tile_X8Y0_S2BEGb;
	wire [15:0] Tile_X8Y0_S4BEG;
	wire [15:0] Tile_X8Y0_SS4BEG;
	wire [3:0] Tile_X9Y0_S1BEG;
	wire [7:0] Tile_X9Y0_S2BEG;
	wire [7:0] Tile_X9Y0_S2BEGb;
	wire [15:0] Tile_X9Y0_S4BEG;
	wire [15:0] Tile_X9Y0_SS4BEG;
	wire [3:0] Tile_X10Y0_S1BEG;
	wire [7:0] Tile_X10Y0_S2BEG;
	wire [7:0] Tile_X10Y0_S2BEGb;
	wire [15:0] Tile_X10Y0_S4BEG;
	wire [15:0] Tile_X10Y0_SS4BEG;
	wire [3:0] Tile_X4Y1_E1BEG;
	wire [7:0] Tile_X4Y1_E2BEG;
	wire [7:0] Tile_X4Y1_E2BEGb;
	wire [15:0] Tile_X4Y1_EE4BEG;
	wire [11:0] Tile_X4Y1_E6BEG;
	wire [3:0] Tile_X5Y1_N1BEG;
	wire [7:0] Tile_X5Y1_N2BEG;
	wire [7:0] Tile_X5Y1_N2BEGb;
	wire [15:0] Tile_X5Y1_N4BEG;
	wire [15:0] Tile_X5Y1_NN4BEG;
	wire [3:0] Tile_X5Y1_E1BEG;
	wire [7:0] Tile_X5Y1_E2BEG;
	wire [7:0] Tile_X5Y1_E2BEGb;
	wire [15:0] Tile_X5Y1_EE4BEG;
	wire [11:0] Tile_X5Y1_E6BEG;
	wire [3:0] Tile_X5Y1_S1BEG;
	wire [7:0] Tile_X5Y1_S2BEG;
	wire [7:0] Tile_X5Y1_S2BEGb;
	wire [15:0] Tile_X5Y1_S4BEG;
	wire [15:0] Tile_X5Y1_SS4BEG;
	wire [17:0] Tile_X5Y1_top2bot;
	wire [3:0] Tile_X5Y1_W1BEG;
	wire [7:0] Tile_X5Y1_W2BEG;
	wire [7:0] Tile_X5Y1_W2BEGb;
	wire [15:0] Tile_X5Y1_WW4BEG;
	wire [11:0] Tile_X5Y1_W6BEG;
	wire [3:0] Tile_X6Y1_N1BEG;
	wire [7:0] Tile_X6Y1_N2BEG;
	wire [7:0] Tile_X6Y1_N2BEGb;
	wire [15:0] Tile_X6Y1_N4BEG;
	wire [15:0] Tile_X6Y1_NN4BEG;
	wire [0:0] Tile_X6Y1_Co;
	wire [3:0] Tile_X6Y1_E1BEG;
	wire [7:0] Tile_X6Y1_E2BEG;
	wire [7:0] Tile_X6Y1_E2BEGb;
	wire [15:0] Tile_X6Y1_EE4BEG;
	wire [11:0] Tile_X6Y1_E6BEG;
	wire [3:0] Tile_X6Y1_S1BEG;
	wire [7:0] Tile_X6Y1_S2BEG;
	wire [7:0] Tile_X6Y1_S2BEGb;
	wire [15:0] Tile_X6Y1_S4BEG;
	wire [15:0] Tile_X6Y1_SS4BEG;
	wire [3:0] Tile_X6Y1_W1BEG;
	wire [7:0] Tile_X6Y1_W2BEG;
	wire [7:0] Tile_X6Y1_W2BEGb;
	wire [15:0] Tile_X6Y1_WW4BEG;
	wire [11:0] Tile_X6Y1_W6BEG;
	wire [3:0] Tile_X7Y1_N1BEG;
	wire [7:0] Tile_X7Y1_N2BEG;
	wire [7:0] Tile_X7Y1_N2BEGb;
	wire [15:0] Tile_X7Y1_N4BEG;
	wire [15:0] Tile_X7Y1_NN4BEG;
	wire [0:0] Tile_X7Y1_Co;
	wire [3:0] Tile_X7Y1_E1BEG;
	wire [7:0] Tile_X7Y1_E2BEG;
	wire [7:0] Tile_X7Y1_E2BEGb;
	wire [15:0] Tile_X7Y1_EE4BEG;
	wire [11:0] Tile_X7Y1_E6BEG;
	wire [3:0] Tile_X7Y1_S1BEG;
	wire [7:0] Tile_X7Y1_S2BEG;
	wire [7:0] Tile_X7Y1_S2BEGb;
	wire [15:0] Tile_X7Y1_S4BEG;
	wire [15:0] Tile_X7Y1_SS4BEG;
	wire [3:0] Tile_X7Y1_W1BEG;
	wire [7:0] Tile_X7Y1_W2BEG;
	wire [7:0] Tile_X7Y1_W2BEGb;
	wire [15:0] Tile_X7Y1_WW4BEG;
	wire [11:0] Tile_X7Y1_W6BEG;
	wire [3:0] Tile_X8Y1_N1BEG;
	wire [7:0] Tile_X8Y1_N2BEG;
	wire [7:0] Tile_X8Y1_N2BEGb;
	wire [15:0] Tile_X8Y1_N4BEG;
	wire [15:0] Tile_X8Y1_NN4BEG;
	wire [0:0] Tile_X8Y1_Co;
	wire [3:0] Tile_X8Y1_E1BEG;
	wire [7:0] Tile_X8Y1_E2BEG;
	wire [7:0] Tile_X8Y1_E2BEGb;
	wire [15:0] Tile_X8Y1_EE4BEG;
	wire [11:0] Tile_X8Y1_E6BEG;
	wire [3:0] Tile_X8Y1_S1BEG;
	wire [7:0] Tile_X8Y1_S2BEG;
	wire [7:0] Tile_X8Y1_S2BEGb;
	wire [15:0] Tile_X8Y1_S4BEG;
	wire [15:0] Tile_X8Y1_SS4BEG;
	wire [3:0] Tile_X8Y1_W1BEG;
	wire [7:0] Tile_X8Y1_W2BEG;
	wire [7:0] Tile_X8Y1_W2BEGb;
	wire [15:0] Tile_X8Y1_WW4BEG;
	wire [11:0] Tile_X8Y1_W6BEG;
	wire [3:0] Tile_X9Y1_N1BEG;
	wire [7:0] Tile_X9Y1_N2BEG;
	wire [7:0] Tile_X9Y1_N2BEGb;
	wire [15:0] Tile_X9Y1_N4BEG;
	wire [15:0] Tile_X9Y1_NN4BEG;
	wire [3:0] Tile_X9Y1_E1BEG;
	wire [7:0] Tile_X9Y1_E2BEG;
	wire [7:0] Tile_X9Y1_E2BEGb;
	wire [15:0] Tile_X9Y1_EE4BEG;
	wire [11:0] Tile_X9Y1_E6BEG;
	wire [3:0] Tile_X9Y1_S1BEG;
	wire [7:0] Tile_X9Y1_S2BEG;
	wire [7:0] Tile_X9Y1_S2BEGb;
	wire [15:0] Tile_X9Y1_S4BEG;
	wire [15:0] Tile_X9Y1_SS4BEG;
	wire [17:0] Tile_X9Y1_top2bot;
	wire [3:0] Tile_X9Y1_W1BEG;
	wire [7:0] Tile_X9Y1_W2BEG;
	wire [7:0] Tile_X9Y1_W2BEGb;
	wire [15:0] Tile_X9Y1_WW4BEG;
	wire [11:0] Tile_X9Y1_W6BEG;
	wire [3:0] Tile_X10Y1_N1BEG;
	wire [7:0] Tile_X10Y1_N2BEG;
	wire [7:0] Tile_X10Y1_N2BEGb;
	wire [15:0] Tile_X10Y1_N4BEG;
	wire [15:0] Tile_X10Y1_NN4BEG;
	wire [0:0] Tile_X10Y1_Co;
	wire [3:0] Tile_X10Y1_E1BEG;
	wire [7:0] Tile_X10Y1_E2BEG;
	wire [7:0] Tile_X10Y1_E2BEGb;
	wire [15:0] Tile_X10Y1_EE4BEG;
	wire [11:0] Tile_X10Y1_E6BEG;
	wire [3:0] Tile_X10Y1_S1BEG;
	wire [7:0] Tile_X10Y1_S2BEG;
	wire [7:0] Tile_X10Y1_S2BEGb;
	wire [15:0] Tile_X10Y1_S4BEG;
	wire [15:0] Tile_X10Y1_SS4BEG;
	wire [3:0] Tile_X10Y1_W1BEG;
	wire [7:0] Tile_X10Y1_W2BEG;
	wire [7:0] Tile_X10Y1_W2BEGb;
	wire [15:0] Tile_X10Y1_WW4BEG;
	wire [11:0] Tile_X10Y1_W6BEG;
	wire [3:0] Tile_X11Y1_W1BEG;
	wire [7:0] Tile_X11Y1_W2BEG;
	wire [7:0] Tile_X11Y1_W2BEGb;
	wire [15:0] Tile_X11Y1_WW4BEG;
	wire [11:0] Tile_X11Y1_W6BEG;
	wire [3:0] Tile_X4Y2_E1BEG;
	wire [7:0] Tile_X4Y2_E2BEG;
	wire [7:0] Tile_X4Y2_E2BEGb;
	wire [15:0] Tile_X4Y2_EE4BEG;
	wire [11:0] Tile_X4Y2_E6BEG;
	wire [3:0] Tile_X5Y2_N1BEG;
	wire [7:0] Tile_X5Y2_N2BEG;
	wire [7:0] Tile_X5Y2_N2BEGb;
	wire [15:0] Tile_X5Y2_N4BEG;
	wire [15:0] Tile_X5Y2_NN4BEG;
	wire [9:0] Tile_X5Y2_bot2top;
	wire [3:0] Tile_X5Y2_E1BEG;
	wire [7:0] Tile_X5Y2_E2BEG;
	wire [7:0] Tile_X5Y2_E2BEGb;
	wire [15:0] Tile_X5Y2_EE4BEG;
	wire [11:0] Tile_X5Y2_E6BEG;
	wire [3:0] Tile_X5Y2_S1BEG;
	wire [7:0] Tile_X5Y2_S2BEG;
	wire [7:0] Tile_X5Y2_S2BEGb;
	wire [15:0] Tile_X5Y2_S4BEG;
	wire [15:0] Tile_X5Y2_SS4BEG;
	wire [3:0] Tile_X5Y2_W1BEG;
	wire [7:0] Tile_X5Y2_W2BEG;
	wire [7:0] Tile_X5Y2_W2BEGb;
	wire [15:0] Tile_X5Y2_WW4BEG;
	wire [11:0] Tile_X5Y2_W6BEG;
	wire [3:0] Tile_X6Y2_N1BEG;
	wire [7:0] Tile_X6Y2_N2BEG;
	wire [7:0] Tile_X6Y2_N2BEGb;
	wire [15:0] Tile_X6Y2_N4BEG;
	wire [15:0] Tile_X6Y2_NN4BEG;
	wire [0:0] Tile_X6Y2_Co;
	wire [3:0] Tile_X6Y2_E1BEG;
	wire [7:0] Tile_X6Y2_E2BEG;
	wire [7:0] Tile_X6Y2_E2BEGb;
	wire [15:0] Tile_X6Y2_EE4BEG;
	wire [11:0] Tile_X6Y2_E6BEG;
	wire [3:0] Tile_X6Y2_S1BEG;
	wire [7:0] Tile_X6Y2_S2BEG;
	wire [7:0] Tile_X6Y2_S2BEGb;
	wire [15:0] Tile_X6Y2_S4BEG;
	wire [15:0] Tile_X6Y2_SS4BEG;
	wire [3:0] Tile_X6Y2_W1BEG;
	wire [7:0] Tile_X6Y2_W2BEG;
	wire [7:0] Tile_X6Y2_W2BEGb;
	wire [15:0] Tile_X6Y2_WW4BEG;
	wire [11:0] Tile_X6Y2_W6BEG;
	wire [3:0] Tile_X7Y2_N1BEG;
	wire [7:0] Tile_X7Y2_N2BEG;
	wire [7:0] Tile_X7Y2_N2BEGb;
	wire [15:0] Tile_X7Y2_N4BEG;
	wire [15:0] Tile_X7Y2_NN4BEG;
	wire [0:0] Tile_X7Y2_Co;
	wire [3:0] Tile_X7Y2_E1BEG;
	wire [7:0] Tile_X7Y2_E2BEG;
	wire [7:0] Tile_X7Y2_E2BEGb;
	wire [15:0] Tile_X7Y2_EE4BEG;
	wire [11:0] Tile_X7Y2_E6BEG;
	wire [3:0] Tile_X7Y2_S1BEG;
	wire [7:0] Tile_X7Y2_S2BEG;
	wire [7:0] Tile_X7Y2_S2BEGb;
	wire [15:0] Tile_X7Y2_S4BEG;
	wire [15:0] Tile_X7Y2_SS4BEG;
	wire [3:0] Tile_X7Y2_W1BEG;
	wire [7:0] Tile_X7Y2_W2BEG;
	wire [7:0] Tile_X7Y2_W2BEGb;
	wire [15:0] Tile_X7Y2_WW4BEG;
	wire [11:0] Tile_X7Y2_W6BEG;
	wire [3:0] Tile_X8Y2_N1BEG;
	wire [7:0] Tile_X8Y2_N2BEG;
	wire [7:0] Tile_X8Y2_N2BEGb;
	wire [15:0] Tile_X8Y2_N4BEG;
	wire [15:0] Tile_X8Y2_NN4BEG;
	wire [0:0] Tile_X8Y2_Co;
	wire [3:0] Tile_X8Y2_E1BEG;
	wire [7:0] Tile_X8Y2_E2BEG;
	wire [7:0] Tile_X8Y2_E2BEGb;
	wire [15:0] Tile_X8Y2_EE4BEG;
	wire [11:0] Tile_X8Y2_E6BEG;
	wire [3:0] Tile_X8Y2_S1BEG;
	wire [7:0] Tile_X8Y2_S2BEG;
	wire [7:0] Tile_X8Y2_S2BEGb;
	wire [15:0] Tile_X8Y2_S4BEG;
	wire [15:0] Tile_X8Y2_SS4BEG;
	wire [3:0] Tile_X8Y2_W1BEG;
	wire [7:0] Tile_X8Y2_W2BEG;
	wire [7:0] Tile_X8Y2_W2BEGb;
	wire [15:0] Tile_X8Y2_WW4BEG;
	wire [11:0] Tile_X8Y2_W6BEG;
	wire [3:0] Tile_X9Y2_N1BEG;
	wire [7:0] Tile_X9Y2_N2BEG;
	wire [7:0] Tile_X9Y2_N2BEGb;
	wire [15:0] Tile_X9Y2_N4BEG;
	wire [15:0] Tile_X9Y2_NN4BEG;
	wire [9:0] Tile_X9Y2_bot2top;
	wire [3:0] Tile_X9Y2_E1BEG;
	wire [7:0] Tile_X9Y2_E2BEG;
	wire [7:0] Tile_X9Y2_E2BEGb;
	wire [15:0] Tile_X9Y2_EE4BEG;
	wire [11:0] Tile_X9Y2_E6BEG;
	wire [3:0] Tile_X9Y2_S1BEG;
	wire [7:0] Tile_X9Y2_S2BEG;
	wire [7:0] Tile_X9Y2_S2BEGb;
	wire [15:0] Tile_X9Y2_S4BEG;
	wire [15:0] Tile_X9Y2_SS4BEG;
	wire [3:0] Tile_X9Y2_W1BEG;
	wire [7:0] Tile_X9Y2_W2BEG;
	wire [7:0] Tile_X9Y2_W2BEGb;
	wire [15:0] Tile_X9Y2_WW4BEG;
	wire [11:0] Tile_X9Y2_W6BEG;
	wire [3:0] Tile_X10Y2_N1BEG;
	wire [7:0] Tile_X10Y2_N2BEG;
	wire [7:0] Tile_X10Y2_N2BEGb;
	wire [15:0] Tile_X10Y2_N4BEG;
	wire [15:0] Tile_X10Y2_NN4BEG;
	wire [0:0] Tile_X10Y2_Co;
	wire [3:0] Tile_X10Y2_E1BEG;
	wire [7:0] Tile_X10Y2_E2BEG;
	wire [7:0] Tile_X10Y2_E2BEGb;
	wire [15:0] Tile_X10Y2_EE4BEG;
	wire [11:0] Tile_X10Y2_E6BEG;
	wire [3:0] Tile_X10Y2_S1BEG;
	wire [7:0] Tile_X10Y2_S2BEG;
	wire [7:0] Tile_X10Y2_S2BEGb;
	wire [15:0] Tile_X10Y2_S4BEG;
	wire [15:0] Tile_X10Y2_SS4BEG;
	wire [3:0] Tile_X10Y2_W1BEG;
	wire [7:0] Tile_X10Y2_W2BEG;
	wire [7:0] Tile_X10Y2_W2BEGb;
	wire [15:0] Tile_X10Y2_WW4BEG;
	wire [11:0] Tile_X10Y2_W6BEG;
	wire [3:0] Tile_X11Y2_W1BEG;
	wire [7:0] Tile_X11Y2_W2BEG;
	wire [7:0] Tile_X11Y2_W2BEGb;
	wire [15:0] Tile_X11Y2_WW4BEG;
	wire [11:0] Tile_X11Y2_W6BEG;
	wire [3:0] Tile_X4Y3_E1BEG;
	wire [7:0] Tile_X4Y3_E2BEG;
	wire [7:0] Tile_X4Y3_E2BEGb;
	wire [15:0] Tile_X4Y3_EE4BEG;
	wire [11:0] Tile_X4Y3_E6BEG;
	wire [3:0] Tile_X5Y3_N1BEG;
	wire [7:0] Tile_X5Y3_N2BEG;
	wire [7:0] Tile_X5Y3_N2BEGb;
	wire [15:0] Tile_X5Y3_N4BEG;
	wire [15:0] Tile_X5Y3_NN4BEG;
	wire [3:0] Tile_X5Y3_E1BEG;
	wire [7:0] Tile_X5Y3_E2BEG;
	wire [7:0] Tile_X5Y3_E2BEGb;
	wire [15:0] Tile_X5Y3_EE4BEG;
	wire [11:0] Tile_X5Y3_E6BEG;
	wire [3:0] Tile_X5Y3_S1BEG;
	wire [7:0] Tile_X5Y3_S2BEG;
	wire [7:0] Tile_X5Y3_S2BEGb;
	wire [15:0] Tile_X5Y3_S4BEG;
	wire [15:0] Tile_X5Y3_SS4BEG;
	wire [17:0] Tile_X5Y3_top2bot;
	wire [3:0] Tile_X5Y3_W1BEG;
	wire [7:0] Tile_X5Y3_W2BEG;
	wire [7:0] Tile_X5Y3_W2BEGb;
	wire [15:0] Tile_X5Y3_WW4BEG;
	wire [11:0] Tile_X5Y3_W6BEG;
	wire [3:0] Tile_X6Y3_N1BEG;
	wire [7:0] Tile_X6Y3_N2BEG;
	wire [7:0] Tile_X6Y3_N2BEGb;
	wire [15:0] Tile_X6Y3_N4BEG;
	wire [15:0] Tile_X6Y3_NN4BEG;
	wire [0:0] Tile_X6Y3_Co;
	wire [3:0] Tile_X6Y3_E1BEG;
	wire [7:0] Tile_X6Y3_E2BEG;
	wire [7:0] Tile_X6Y3_E2BEGb;
	wire [15:0] Tile_X6Y3_EE4BEG;
	wire [11:0] Tile_X6Y3_E6BEG;
	wire [3:0] Tile_X6Y3_S1BEG;
	wire [7:0] Tile_X6Y3_S2BEG;
	wire [7:0] Tile_X6Y3_S2BEGb;
	wire [15:0] Tile_X6Y3_S4BEG;
	wire [15:0] Tile_X6Y3_SS4BEG;
	wire [3:0] Tile_X6Y3_W1BEG;
	wire [7:0] Tile_X6Y3_W2BEG;
	wire [7:0] Tile_X6Y3_W2BEGb;
	wire [15:0] Tile_X6Y3_WW4BEG;
	wire [11:0] Tile_X6Y3_W6BEG;
	wire [3:0] Tile_X7Y3_N1BEG;
	wire [7:0] Tile_X7Y3_N2BEG;
	wire [7:0] Tile_X7Y3_N2BEGb;
	wire [15:0] Tile_X7Y3_N4BEG;
	wire [15:0] Tile_X7Y3_NN4BEG;
	wire [0:0] Tile_X7Y3_Co;
	wire [3:0] Tile_X7Y3_E1BEG;
	wire [7:0] Tile_X7Y3_E2BEG;
	wire [7:0] Tile_X7Y3_E2BEGb;
	wire [15:0] Tile_X7Y3_EE4BEG;
	wire [11:0] Tile_X7Y3_E6BEG;
	wire [3:0] Tile_X7Y3_S1BEG;
	wire [7:0] Tile_X7Y3_S2BEG;
	wire [7:0] Tile_X7Y3_S2BEGb;
	wire [15:0] Tile_X7Y3_S4BEG;
	wire [15:0] Tile_X7Y3_SS4BEG;
	wire [3:0] Tile_X7Y3_W1BEG;
	wire [7:0] Tile_X7Y3_W2BEG;
	wire [7:0] Tile_X7Y3_W2BEGb;
	wire [15:0] Tile_X7Y3_WW4BEG;
	wire [11:0] Tile_X7Y3_W6BEG;
	wire [3:0] Tile_X8Y3_N1BEG;
	wire [7:0] Tile_X8Y3_N2BEG;
	wire [7:0] Tile_X8Y3_N2BEGb;
	wire [15:0] Tile_X8Y3_N4BEG;
	wire [15:0] Tile_X8Y3_NN4BEG;
	wire [0:0] Tile_X8Y3_Co;
	wire [3:0] Tile_X8Y3_E1BEG;
	wire [7:0] Tile_X8Y3_E2BEG;
	wire [7:0] Tile_X8Y3_E2BEGb;
	wire [15:0] Tile_X8Y3_EE4BEG;
	wire [11:0] Tile_X8Y3_E6BEG;
	wire [3:0] Tile_X8Y3_S1BEG;
	wire [7:0] Tile_X8Y3_S2BEG;
	wire [7:0] Tile_X8Y3_S2BEGb;
	wire [15:0] Tile_X8Y3_S4BEG;
	wire [15:0] Tile_X8Y3_SS4BEG;
	wire [3:0] Tile_X8Y3_W1BEG;
	wire [7:0] Tile_X8Y3_W2BEG;
	wire [7:0] Tile_X8Y3_W2BEGb;
	wire [15:0] Tile_X8Y3_WW4BEG;
	wire [11:0] Tile_X8Y3_W6BEG;
	wire [3:0] Tile_X9Y3_N1BEG;
	wire [7:0] Tile_X9Y3_N2BEG;
	wire [7:0] Tile_X9Y3_N2BEGb;
	wire [15:0] Tile_X9Y3_N4BEG;
	wire [15:0] Tile_X9Y3_NN4BEG;
	wire [3:0] Tile_X9Y3_E1BEG;
	wire [7:0] Tile_X9Y3_E2BEG;
	wire [7:0] Tile_X9Y3_E2BEGb;
	wire [15:0] Tile_X9Y3_EE4BEG;
	wire [11:0] Tile_X9Y3_E6BEG;
	wire [3:0] Tile_X9Y3_S1BEG;
	wire [7:0] Tile_X9Y3_S2BEG;
	wire [7:0] Tile_X9Y3_S2BEGb;
	wire [15:0] Tile_X9Y3_S4BEG;
	wire [15:0] Tile_X9Y3_SS4BEG;
	wire [17:0] Tile_X9Y3_top2bot;
	wire [3:0] Tile_X9Y3_W1BEG;
	wire [7:0] Tile_X9Y3_W2BEG;
	wire [7:0] Tile_X9Y3_W2BEGb;
	wire [15:0] Tile_X9Y3_WW4BEG;
	wire [11:0] Tile_X9Y3_W6BEG;
	wire [3:0] Tile_X10Y3_N1BEG;
	wire [7:0] Tile_X10Y3_N2BEG;
	wire [7:0] Tile_X10Y3_N2BEGb;
	wire [15:0] Tile_X10Y3_N4BEG;
	wire [15:0] Tile_X10Y3_NN4BEG;
	wire [0:0] Tile_X10Y3_Co;
	wire [3:0] Tile_X10Y3_E1BEG;
	wire [7:0] Tile_X10Y3_E2BEG;
	wire [7:0] Tile_X10Y3_E2BEGb;
	wire [15:0] Tile_X10Y3_EE4BEG;
	wire [11:0] Tile_X10Y3_E6BEG;
	wire [3:0] Tile_X10Y3_S1BEG;
	wire [7:0] Tile_X10Y3_S2BEG;
	wire [7:0] Tile_X10Y3_S2BEGb;
	wire [15:0] Tile_X10Y3_S4BEG;
	wire [15:0] Tile_X10Y3_SS4BEG;
	wire [3:0] Tile_X10Y3_W1BEG;
	wire [7:0] Tile_X10Y3_W2BEG;
	wire [7:0] Tile_X10Y3_W2BEGb;
	wire [15:0] Tile_X10Y3_WW4BEG;
	wire [11:0] Tile_X10Y3_W6BEG;
	wire [3:0] Tile_X11Y3_W1BEG;
	wire [7:0] Tile_X11Y3_W2BEG;
	wire [7:0] Tile_X11Y3_W2BEGb;
	wire [15:0] Tile_X11Y3_WW4BEG;
	wire [11:0] Tile_X11Y3_W6BEG;
	wire [3:0] Tile_X4Y4_E1BEG;
	wire [7:0] Tile_X4Y4_E2BEG;
	wire [7:0] Tile_X4Y4_E2BEGb;
	wire [15:0] Tile_X4Y4_EE4BEG;
	wire [11:0] Tile_X4Y4_E6BEG;
	wire [3:0] Tile_X5Y4_N1BEG;
	wire [7:0] Tile_X5Y4_N2BEG;
	wire [7:0] Tile_X5Y4_N2BEGb;
	wire [15:0] Tile_X5Y4_N4BEG;
	wire [15:0] Tile_X5Y4_NN4BEG;
	wire [9:0] Tile_X5Y4_bot2top;
	wire [3:0] Tile_X5Y4_E1BEG;
	wire [7:0] Tile_X5Y4_E2BEG;
	wire [7:0] Tile_X5Y4_E2BEGb;
	wire [15:0] Tile_X5Y4_EE4BEG;
	wire [11:0] Tile_X5Y4_E6BEG;
	wire [3:0] Tile_X5Y4_S1BEG;
	wire [7:0] Tile_X5Y4_S2BEG;
	wire [7:0] Tile_X5Y4_S2BEGb;
	wire [15:0] Tile_X5Y4_S4BEG;
	wire [15:0] Tile_X5Y4_SS4BEG;
	wire [3:0] Tile_X5Y4_W1BEG;
	wire [7:0] Tile_X5Y4_W2BEG;
	wire [7:0] Tile_X5Y4_W2BEGb;
	wire [15:0] Tile_X5Y4_WW4BEG;
	wire [11:0] Tile_X5Y4_W6BEG;
	wire [3:0] Tile_X6Y4_N1BEG;
	wire [7:0] Tile_X6Y4_N2BEG;
	wire [7:0] Tile_X6Y4_N2BEGb;
	wire [15:0] Tile_X6Y4_N4BEG;
	wire [15:0] Tile_X6Y4_NN4BEG;
	wire [0:0] Tile_X6Y4_Co;
	wire [3:0] Tile_X6Y4_E1BEG;
	wire [7:0] Tile_X6Y4_E2BEG;
	wire [7:0] Tile_X6Y4_E2BEGb;
	wire [15:0] Tile_X6Y4_EE4BEG;
	wire [11:0] Tile_X6Y4_E6BEG;
	wire [3:0] Tile_X6Y4_S1BEG;
	wire [7:0] Tile_X6Y4_S2BEG;
	wire [7:0] Tile_X6Y4_S2BEGb;
	wire [15:0] Tile_X6Y4_S4BEG;
	wire [15:0] Tile_X6Y4_SS4BEG;
	wire [3:0] Tile_X6Y4_W1BEG;
	wire [7:0] Tile_X6Y4_W2BEG;
	wire [7:0] Tile_X6Y4_W2BEGb;
	wire [15:0] Tile_X6Y4_WW4BEG;
	wire [11:0] Tile_X6Y4_W6BEG;
	wire [3:0] Tile_X7Y4_N1BEG;
	wire [7:0] Tile_X7Y4_N2BEG;
	wire [7:0] Tile_X7Y4_N2BEGb;
	wire [15:0] Tile_X7Y4_N4BEG;
	wire [15:0] Tile_X7Y4_NN4BEG;
	wire [0:0] Tile_X7Y4_Co;
	wire [3:0] Tile_X7Y4_E1BEG;
	wire [7:0] Tile_X7Y4_E2BEG;
	wire [7:0] Tile_X7Y4_E2BEGb;
	wire [15:0] Tile_X7Y4_EE4BEG;
	wire [11:0] Tile_X7Y4_E6BEG;
	wire [3:0] Tile_X7Y4_S1BEG;
	wire [7:0] Tile_X7Y4_S2BEG;
	wire [7:0] Tile_X7Y4_S2BEGb;
	wire [15:0] Tile_X7Y4_S4BEG;
	wire [15:0] Tile_X7Y4_SS4BEG;
	wire [3:0] Tile_X7Y4_W1BEG;
	wire [7:0] Tile_X7Y4_W2BEG;
	wire [7:0] Tile_X7Y4_W2BEGb;
	wire [15:0] Tile_X7Y4_WW4BEG;
	wire [11:0] Tile_X7Y4_W6BEG;
	wire [3:0] Tile_X8Y4_N1BEG;
	wire [7:0] Tile_X8Y4_N2BEG;
	wire [7:0] Tile_X8Y4_N2BEGb;
	wire [15:0] Tile_X8Y4_N4BEG;
	wire [15:0] Tile_X8Y4_NN4BEG;
	wire [0:0] Tile_X8Y4_Co;
	wire [3:0] Tile_X8Y4_E1BEG;
	wire [7:0] Tile_X8Y4_E2BEG;
	wire [7:0] Tile_X8Y4_E2BEGb;
	wire [15:0] Tile_X8Y4_EE4BEG;
	wire [11:0] Tile_X8Y4_E6BEG;
	wire [3:0] Tile_X8Y4_S1BEG;
	wire [7:0] Tile_X8Y4_S2BEG;
	wire [7:0] Tile_X8Y4_S2BEGb;
	wire [15:0] Tile_X8Y4_S4BEG;
	wire [15:0] Tile_X8Y4_SS4BEG;
	wire [3:0] Tile_X8Y4_W1BEG;
	wire [7:0] Tile_X8Y4_W2BEG;
	wire [7:0] Tile_X8Y4_W2BEGb;
	wire [15:0] Tile_X8Y4_WW4BEG;
	wire [11:0] Tile_X8Y4_W6BEG;
	wire [3:0] Tile_X9Y4_N1BEG;
	wire [7:0] Tile_X9Y4_N2BEG;
	wire [7:0] Tile_X9Y4_N2BEGb;
	wire [15:0] Tile_X9Y4_N4BEG;
	wire [15:0] Tile_X9Y4_NN4BEG;
	wire [9:0] Tile_X9Y4_bot2top;
	wire [3:0] Tile_X9Y4_E1BEG;
	wire [7:0] Tile_X9Y4_E2BEG;
	wire [7:0] Tile_X9Y4_E2BEGb;
	wire [15:0] Tile_X9Y4_EE4BEG;
	wire [11:0] Tile_X9Y4_E6BEG;
	wire [3:0] Tile_X9Y4_S1BEG;
	wire [7:0] Tile_X9Y4_S2BEG;
	wire [7:0] Tile_X9Y4_S2BEGb;
	wire [15:0] Tile_X9Y4_S4BEG;
	wire [15:0] Tile_X9Y4_SS4BEG;
	wire [3:0] Tile_X9Y4_W1BEG;
	wire [7:0] Tile_X9Y4_W2BEG;
	wire [7:0] Tile_X9Y4_W2BEGb;
	wire [15:0] Tile_X9Y4_WW4BEG;
	wire [11:0] Tile_X9Y4_W6BEG;
	wire [3:0] Tile_X10Y4_N1BEG;
	wire [7:0] Tile_X10Y4_N2BEG;
	wire [7:0] Tile_X10Y4_N2BEGb;
	wire [15:0] Tile_X10Y4_N4BEG;
	wire [15:0] Tile_X10Y4_NN4BEG;
	wire [0:0] Tile_X10Y4_Co;
	wire [3:0] Tile_X10Y4_E1BEG;
	wire [7:0] Tile_X10Y4_E2BEG;
	wire [7:0] Tile_X10Y4_E2BEGb;
	wire [15:0] Tile_X10Y4_EE4BEG;
	wire [11:0] Tile_X10Y4_E6BEG;
	wire [3:0] Tile_X10Y4_S1BEG;
	wire [7:0] Tile_X10Y4_S2BEG;
	wire [7:0] Tile_X10Y4_S2BEGb;
	wire [15:0] Tile_X10Y4_S4BEG;
	wire [15:0] Tile_X10Y4_SS4BEG;
	wire [3:0] Tile_X10Y4_W1BEG;
	wire [7:0] Tile_X10Y4_W2BEG;
	wire [7:0] Tile_X10Y4_W2BEGb;
	wire [15:0] Tile_X10Y4_WW4BEG;
	wire [11:0] Tile_X10Y4_W6BEG;
	wire [3:0] Tile_X11Y4_W1BEG;
	wire [7:0] Tile_X11Y4_W2BEG;
	wire [7:0] Tile_X11Y4_W2BEGb;
	wire [15:0] Tile_X11Y4_WW4BEG;
	wire [11:0] Tile_X11Y4_W6BEG;
	wire [3:0] Tile_X4Y5_E1BEG;
	wire [7:0] Tile_X4Y5_E2BEG;
	wire [7:0] Tile_X4Y5_E2BEGb;
	wire [15:0] Tile_X4Y5_EE4BEG;
	wire [11:0] Tile_X4Y5_E6BEG;
	wire [3:0] Tile_X5Y5_N1BEG;
	wire [7:0] Tile_X5Y5_N2BEG;
	wire [7:0] Tile_X5Y5_N2BEGb;
	wire [15:0] Tile_X5Y5_N4BEG;
	wire [15:0] Tile_X5Y5_NN4BEG;
	wire [3:0] Tile_X5Y5_E1BEG;
	wire [7:0] Tile_X5Y5_E2BEG;
	wire [7:0] Tile_X5Y5_E2BEGb;
	wire [15:0] Tile_X5Y5_EE4BEG;
	wire [11:0] Tile_X5Y5_E6BEG;
	wire [3:0] Tile_X5Y5_S1BEG;
	wire [7:0] Tile_X5Y5_S2BEG;
	wire [7:0] Tile_X5Y5_S2BEGb;
	wire [15:0] Tile_X5Y5_S4BEG;
	wire [15:0] Tile_X5Y5_SS4BEG;
	wire [17:0] Tile_X5Y5_top2bot;
	wire [3:0] Tile_X5Y5_W1BEG;
	wire [7:0] Tile_X5Y5_W2BEG;
	wire [7:0] Tile_X5Y5_W2BEGb;
	wire [15:0] Tile_X5Y5_WW4BEG;
	wire [11:0] Tile_X5Y5_W6BEG;
	wire [3:0] Tile_X6Y5_N1BEG;
	wire [7:0] Tile_X6Y5_N2BEG;
	wire [7:0] Tile_X6Y5_N2BEGb;
	wire [15:0] Tile_X6Y5_N4BEG;
	wire [15:0] Tile_X6Y5_NN4BEG;
	wire [0:0] Tile_X6Y5_Co;
	wire [3:0] Tile_X6Y5_E1BEG;
	wire [7:0] Tile_X6Y5_E2BEG;
	wire [7:0] Tile_X6Y5_E2BEGb;
	wire [15:0] Tile_X6Y5_EE4BEG;
	wire [11:0] Tile_X6Y5_E6BEG;
	wire [3:0] Tile_X6Y5_S1BEG;
	wire [7:0] Tile_X6Y5_S2BEG;
	wire [7:0] Tile_X6Y5_S2BEGb;
	wire [15:0] Tile_X6Y5_S4BEG;
	wire [15:0] Tile_X6Y5_SS4BEG;
	wire [3:0] Tile_X6Y5_W1BEG;
	wire [7:0] Tile_X6Y5_W2BEG;
	wire [7:0] Tile_X6Y5_W2BEGb;
	wire [15:0] Tile_X6Y5_WW4BEG;
	wire [11:0] Tile_X6Y5_W6BEG;
	wire [3:0] Tile_X7Y5_N1BEG;
	wire [7:0] Tile_X7Y5_N2BEG;
	wire [7:0] Tile_X7Y5_N2BEGb;
	wire [15:0] Tile_X7Y5_N4BEG;
	wire [15:0] Tile_X7Y5_NN4BEG;
	wire [0:0] Tile_X7Y5_Co;
	wire [3:0] Tile_X7Y5_E1BEG;
	wire [7:0] Tile_X7Y5_E2BEG;
	wire [7:0] Tile_X7Y5_E2BEGb;
	wire [15:0] Tile_X7Y5_EE4BEG;
	wire [11:0] Tile_X7Y5_E6BEG;
	wire [3:0] Tile_X7Y5_S1BEG;
	wire [7:0] Tile_X7Y5_S2BEG;
	wire [7:0] Tile_X7Y5_S2BEGb;
	wire [15:0] Tile_X7Y5_S4BEG;
	wire [15:0] Tile_X7Y5_SS4BEG;
	wire [3:0] Tile_X7Y5_W1BEG;
	wire [7:0] Tile_X7Y5_W2BEG;
	wire [7:0] Tile_X7Y5_W2BEGb;
	wire [15:0] Tile_X7Y5_WW4BEG;
	wire [11:0] Tile_X7Y5_W6BEG;
	wire [3:0] Tile_X8Y5_N1BEG;
	wire [7:0] Tile_X8Y5_N2BEG;
	wire [7:0] Tile_X8Y5_N2BEGb;
	wire [15:0] Tile_X8Y5_N4BEG;
	wire [15:0] Tile_X8Y5_NN4BEG;
	wire [0:0] Tile_X8Y5_Co;
	wire [3:0] Tile_X8Y5_E1BEG;
	wire [7:0] Tile_X8Y5_E2BEG;
	wire [7:0] Tile_X8Y5_E2BEGb;
	wire [15:0] Tile_X8Y5_EE4BEG;
	wire [11:0] Tile_X8Y5_E6BEG;
	wire [3:0] Tile_X8Y5_S1BEG;
	wire [7:0] Tile_X8Y5_S2BEG;
	wire [7:0] Tile_X8Y5_S2BEGb;
	wire [15:0] Tile_X8Y5_S4BEG;
	wire [15:0] Tile_X8Y5_SS4BEG;
	wire [3:0] Tile_X8Y5_W1BEG;
	wire [7:0] Tile_X8Y5_W2BEG;
	wire [7:0] Tile_X8Y5_W2BEGb;
	wire [15:0] Tile_X8Y5_WW4BEG;
	wire [11:0] Tile_X8Y5_W6BEG;
	wire [3:0] Tile_X9Y5_N1BEG;
	wire [7:0] Tile_X9Y5_N2BEG;
	wire [7:0] Tile_X9Y5_N2BEGb;
	wire [15:0] Tile_X9Y5_N4BEG;
	wire [15:0] Tile_X9Y5_NN4BEG;
	wire [3:0] Tile_X9Y5_E1BEG;
	wire [7:0] Tile_X9Y5_E2BEG;
	wire [7:0] Tile_X9Y5_E2BEGb;
	wire [15:0] Tile_X9Y5_EE4BEG;
	wire [11:0] Tile_X9Y5_E6BEG;
	wire [3:0] Tile_X9Y5_S1BEG;
	wire [7:0] Tile_X9Y5_S2BEG;
	wire [7:0] Tile_X9Y5_S2BEGb;
	wire [15:0] Tile_X9Y5_S4BEG;
	wire [15:0] Tile_X9Y5_SS4BEG;
	wire [17:0] Tile_X9Y5_top2bot;
	wire [3:0] Tile_X9Y5_W1BEG;
	wire [7:0] Tile_X9Y5_W2BEG;
	wire [7:0] Tile_X9Y5_W2BEGb;
	wire [15:0] Tile_X9Y5_WW4BEG;
	wire [11:0] Tile_X9Y5_W6BEG;
	wire [3:0] Tile_X10Y5_N1BEG;
	wire [7:0] Tile_X10Y5_N2BEG;
	wire [7:0] Tile_X10Y5_N2BEGb;
	wire [15:0] Tile_X10Y5_N4BEG;
	wire [15:0] Tile_X10Y5_NN4BEG;
	wire [0:0] Tile_X10Y5_Co;
	wire [3:0] Tile_X10Y5_E1BEG;
	wire [7:0] Tile_X10Y5_E2BEG;
	wire [7:0] Tile_X10Y5_E2BEGb;
	wire [15:0] Tile_X10Y5_EE4BEG;
	wire [11:0] Tile_X10Y5_E6BEG;
	wire [3:0] Tile_X10Y5_S1BEG;
	wire [7:0] Tile_X10Y5_S2BEG;
	wire [7:0] Tile_X10Y5_S2BEGb;
	wire [15:0] Tile_X10Y5_S4BEG;
	wire [15:0] Tile_X10Y5_SS4BEG;
	wire [3:0] Tile_X10Y5_W1BEG;
	wire [7:0] Tile_X10Y5_W2BEG;
	wire [7:0] Tile_X10Y5_W2BEGb;
	wire [15:0] Tile_X10Y5_WW4BEG;
	wire [11:0] Tile_X10Y5_W6BEG;
	wire [3:0] Tile_X11Y5_W1BEG;
	wire [7:0] Tile_X11Y5_W2BEG;
	wire [7:0] Tile_X11Y5_W2BEGb;
	wire [15:0] Tile_X11Y5_WW4BEG;
	wire [11:0] Tile_X11Y5_W6BEG;
	wire [3:0] Tile_X4Y6_E1BEG;
	wire [7:0] Tile_X4Y6_E2BEG;
	wire [7:0] Tile_X4Y6_E2BEGb;
	wire [15:0] Tile_X4Y6_EE4BEG;
	wire [11:0] Tile_X4Y6_E6BEG;
	wire [3:0] Tile_X5Y6_N1BEG;
	wire [7:0] Tile_X5Y6_N2BEG;
	wire [7:0] Tile_X5Y6_N2BEGb;
	wire [15:0] Tile_X5Y6_N4BEG;
	wire [15:0] Tile_X5Y6_NN4BEG;
	wire [9:0] Tile_X5Y6_bot2top;
	wire [3:0] Tile_X5Y6_E1BEG;
	wire [7:0] Tile_X5Y6_E2BEG;
	wire [7:0] Tile_X5Y6_E2BEGb;
	wire [15:0] Tile_X5Y6_EE4BEG;
	wire [11:0] Tile_X5Y6_E6BEG;
	wire [3:0] Tile_X5Y6_S1BEG;
	wire [7:0] Tile_X5Y6_S2BEG;
	wire [7:0] Tile_X5Y6_S2BEGb;
	wire [15:0] Tile_X5Y6_S4BEG;
	wire [15:0] Tile_X5Y6_SS4BEG;
	wire [3:0] Tile_X5Y6_W1BEG;
	wire [7:0] Tile_X5Y6_W2BEG;
	wire [7:0] Tile_X5Y6_W2BEGb;
	wire [15:0] Tile_X5Y6_WW4BEG;
	wire [11:0] Tile_X5Y6_W6BEG;
	wire [3:0] Tile_X6Y6_N1BEG;
	wire [7:0] Tile_X6Y6_N2BEG;
	wire [7:0] Tile_X6Y6_N2BEGb;
	wire [15:0] Tile_X6Y6_N4BEG;
	wire [15:0] Tile_X6Y6_NN4BEG;
	wire [0:0] Tile_X6Y6_Co;
	wire [3:0] Tile_X6Y6_E1BEG;
	wire [7:0] Tile_X6Y6_E2BEG;
	wire [7:0] Tile_X6Y6_E2BEGb;
	wire [15:0] Tile_X6Y6_EE4BEG;
	wire [11:0] Tile_X6Y6_E6BEG;
	wire [3:0] Tile_X6Y6_S1BEG;
	wire [7:0] Tile_X6Y6_S2BEG;
	wire [7:0] Tile_X6Y6_S2BEGb;
	wire [15:0] Tile_X6Y6_S4BEG;
	wire [15:0] Tile_X6Y6_SS4BEG;
	wire [3:0] Tile_X6Y6_W1BEG;
	wire [7:0] Tile_X6Y6_W2BEG;
	wire [7:0] Tile_X6Y6_W2BEGb;
	wire [15:0] Tile_X6Y6_WW4BEG;
	wire [11:0] Tile_X6Y6_W6BEG;
	wire [3:0] Tile_X7Y6_N1BEG;
	wire [7:0] Tile_X7Y6_N2BEG;
	wire [7:0] Tile_X7Y6_N2BEGb;
	wire [15:0] Tile_X7Y6_N4BEG;
	wire [15:0] Tile_X7Y6_NN4BEG;
	wire [0:0] Tile_X7Y6_Co;
	wire [3:0] Tile_X7Y6_E1BEG;
	wire [7:0] Tile_X7Y6_E2BEG;
	wire [7:0] Tile_X7Y6_E2BEGb;
	wire [15:0] Tile_X7Y6_EE4BEG;
	wire [11:0] Tile_X7Y6_E6BEG;
	wire [3:0] Tile_X7Y6_S1BEG;
	wire [7:0] Tile_X7Y6_S2BEG;
	wire [7:0] Tile_X7Y6_S2BEGb;
	wire [15:0] Tile_X7Y6_S4BEG;
	wire [15:0] Tile_X7Y6_SS4BEG;
	wire [3:0] Tile_X7Y6_W1BEG;
	wire [7:0] Tile_X7Y6_W2BEG;
	wire [7:0] Tile_X7Y6_W2BEGb;
	wire [15:0] Tile_X7Y6_WW4BEG;
	wire [11:0] Tile_X7Y6_W6BEG;
	wire [3:0] Tile_X8Y6_N1BEG;
	wire [7:0] Tile_X8Y6_N2BEG;
	wire [7:0] Tile_X8Y6_N2BEGb;
	wire [15:0] Tile_X8Y6_N4BEG;
	wire [15:0] Tile_X8Y6_NN4BEG;
	wire [0:0] Tile_X8Y6_Co;
	wire [3:0] Tile_X8Y6_E1BEG;
	wire [7:0] Tile_X8Y6_E2BEG;
	wire [7:0] Tile_X8Y6_E2BEGb;
	wire [15:0] Tile_X8Y6_EE4BEG;
	wire [11:0] Tile_X8Y6_E6BEG;
	wire [3:0] Tile_X8Y6_S1BEG;
	wire [7:0] Tile_X8Y6_S2BEG;
	wire [7:0] Tile_X8Y6_S2BEGb;
	wire [15:0] Tile_X8Y6_S4BEG;
	wire [15:0] Tile_X8Y6_SS4BEG;
	wire [3:0] Tile_X8Y6_W1BEG;
	wire [7:0] Tile_X8Y6_W2BEG;
	wire [7:0] Tile_X8Y6_W2BEGb;
	wire [15:0] Tile_X8Y6_WW4BEG;
	wire [11:0] Tile_X8Y6_W6BEG;
	wire [3:0] Tile_X9Y6_N1BEG;
	wire [7:0] Tile_X9Y6_N2BEG;
	wire [7:0] Tile_X9Y6_N2BEGb;
	wire [15:0] Tile_X9Y6_N4BEG;
	wire [15:0] Tile_X9Y6_NN4BEG;
	wire [9:0] Tile_X9Y6_bot2top;
	wire [3:0] Tile_X9Y6_E1BEG;
	wire [7:0] Tile_X9Y6_E2BEG;
	wire [7:0] Tile_X9Y6_E2BEGb;
	wire [15:0] Tile_X9Y6_EE4BEG;
	wire [11:0] Tile_X9Y6_E6BEG;
	wire [3:0] Tile_X9Y6_S1BEG;
	wire [7:0] Tile_X9Y6_S2BEG;
	wire [7:0] Tile_X9Y6_S2BEGb;
	wire [15:0] Tile_X9Y6_S4BEG;
	wire [15:0] Tile_X9Y6_SS4BEG;
	wire [3:0] Tile_X9Y6_W1BEG;
	wire [7:0] Tile_X9Y6_W2BEG;
	wire [7:0] Tile_X9Y6_W2BEGb;
	wire [15:0] Tile_X9Y6_WW4BEG;
	wire [11:0] Tile_X9Y6_W6BEG;
	wire [3:0] Tile_X10Y6_N1BEG;
	wire [7:0] Tile_X10Y6_N2BEG;
	wire [7:0] Tile_X10Y6_N2BEGb;
	wire [15:0] Tile_X10Y6_N4BEG;
	wire [15:0] Tile_X10Y6_NN4BEG;
	wire [0:0] Tile_X10Y6_Co;
	wire [3:0] Tile_X10Y6_E1BEG;
	wire [7:0] Tile_X10Y6_E2BEG;
	wire [7:0] Tile_X10Y6_E2BEGb;
	wire [15:0] Tile_X10Y6_EE4BEG;
	wire [11:0] Tile_X10Y6_E6BEG;
	wire [3:0] Tile_X10Y6_S1BEG;
	wire [7:0] Tile_X10Y6_S2BEG;
	wire [7:0] Tile_X10Y6_S2BEGb;
	wire [15:0] Tile_X10Y6_S4BEG;
	wire [15:0] Tile_X10Y6_SS4BEG;
	wire [3:0] Tile_X10Y6_W1BEG;
	wire [7:0] Tile_X10Y6_W2BEG;
	wire [7:0] Tile_X10Y6_W2BEGb;
	wire [15:0] Tile_X10Y6_WW4BEG;
	wire [11:0] Tile_X10Y6_W6BEG;
	wire [3:0] Tile_X11Y6_W1BEG;
	wire [7:0] Tile_X11Y6_W2BEG;
	wire [7:0] Tile_X11Y6_W2BEGb;
	wire [15:0] Tile_X11Y6_WW4BEG;
	wire [11:0] Tile_X11Y6_W6BEG;
	wire [3:0] Tile_X4Y7_E1BEG;
	wire [7:0] Tile_X4Y7_E2BEG;
	wire [7:0] Tile_X4Y7_E2BEGb;
	wire [15:0] Tile_X4Y7_EE4BEG;
	wire [11:0] Tile_X4Y7_E6BEG;
	wire [3:0] Tile_X5Y7_N1BEG;
	wire [7:0] Tile_X5Y7_N2BEG;
	wire [7:0] Tile_X5Y7_N2BEGb;
	wire [15:0] Tile_X5Y7_N4BEG;
	wire [15:0] Tile_X5Y7_NN4BEG;
	wire [3:0] Tile_X5Y7_E1BEG;
	wire [7:0] Tile_X5Y7_E2BEG;
	wire [7:0] Tile_X5Y7_E2BEGb;
	wire [15:0] Tile_X5Y7_EE4BEG;
	wire [11:0] Tile_X5Y7_E6BEG;
	wire [3:0] Tile_X5Y7_S1BEG;
	wire [7:0] Tile_X5Y7_S2BEG;
	wire [7:0] Tile_X5Y7_S2BEGb;
	wire [15:0] Tile_X5Y7_S4BEG;
	wire [15:0] Tile_X5Y7_SS4BEG;
	wire [17:0] Tile_X5Y7_top2bot;
	wire [3:0] Tile_X5Y7_W1BEG;
	wire [7:0] Tile_X5Y7_W2BEG;
	wire [7:0] Tile_X5Y7_W2BEGb;
	wire [15:0] Tile_X5Y7_WW4BEG;
	wire [11:0] Tile_X5Y7_W6BEG;
	wire [3:0] Tile_X6Y7_N1BEG;
	wire [7:0] Tile_X6Y7_N2BEG;
	wire [7:0] Tile_X6Y7_N2BEGb;
	wire [15:0] Tile_X6Y7_N4BEG;
	wire [15:0] Tile_X6Y7_NN4BEG;
	wire [0:0] Tile_X6Y7_Co;
	wire [3:0] Tile_X6Y7_E1BEG;
	wire [7:0] Tile_X6Y7_E2BEG;
	wire [7:0] Tile_X6Y7_E2BEGb;
	wire [15:0] Tile_X6Y7_EE4BEG;
	wire [11:0] Tile_X6Y7_E6BEG;
	wire [3:0] Tile_X6Y7_S1BEG;
	wire [7:0] Tile_X6Y7_S2BEG;
	wire [7:0] Tile_X6Y7_S2BEGb;
	wire [15:0] Tile_X6Y7_S4BEG;
	wire [15:0] Tile_X6Y7_SS4BEG;
	wire [3:0] Tile_X6Y7_W1BEG;
	wire [7:0] Tile_X6Y7_W2BEG;
	wire [7:0] Tile_X6Y7_W2BEGb;
	wire [15:0] Tile_X6Y7_WW4BEG;
	wire [11:0] Tile_X6Y7_W6BEG;
	wire [3:0] Tile_X7Y7_N1BEG;
	wire [7:0] Tile_X7Y7_N2BEG;
	wire [7:0] Tile_X7Y7_N2BEGb;
	wire [15:0] Tile_X7Y7_N4BEG;
	wire [15:0] Tile_X7Y7_NN4BEG;
	wire [0:0] Tile_X7Y7_Co;
	wire [3:0] Tile_X7Y7_E1BEG;
	wire [7:0] Tile_X7Y7_E2BEG;
	wire [7:0] Tile_X7Y7_E2BEGb;
	wire [15:0] Tile_X7Y7_EE4BEG;
	wire [11:0] Tile_X7Y7_E6BEG;
	wire [3:0] Tile_X7Y7_S1BEG;
	wire [7:0] Tile_X7Y7_S2BEG;
	wire [7:0] Tile_X7Y7_S2BEGb;
	wire [15:0] Tile_X7Y7_S4BEG;
	wire [15:0] Tile_X7Y7_SS4BEG;
	wire [3:0] Tile_X7Y7_W1BEG;
	wire [7:0] Tile_X7Y7_W2BEG;
	wire [7:0] Tile_X7Y7_W2BEGb;
	wire [15:0] Tile_X7Y7_WW4BEG;
	wire [11:0] Tile_X7Y7_W6BEG;
	wire [3:0] Tile_X8Y7_N1BEG;
	wire [7:0] Tile_X8Y7_N2BEG;
	wire [7:0] Tile_X8Y7_N2BEGb;
	wire [15:0] Tile_X8Y7_N4BEG;
	wire [15:0] Tile_X8Y7_NN4BEG;
	wire [0:0] Tile_X8Y7_Co;
	wire [3:0] Tile_X8Y7_E1BEG;
	wire [7:0] Tile_X8Y7_E2BEG;
	wire [7:0] Tile_X8Y7_E2BEGb;
	wire [15:0] Tile_X8Y7_EE4BEG;
	wire [11:0] Tile_X8Y7_E6BEG;
	wire [3:0] Tile_X8Y7_S1BEG;
	wire [7:0] Tile_X8Y7_S2BEG;
	wire [7:0] Tile_X8Y7_S2BEGb;
	wire [15:0] Tile_X8Y7_S4BEG;
	wire [15:0] Tile_X8Y7_SS4BEG;
	wire [3:0] Tile_X8Y7_W1BEG;
	wire [7:0] Tile_X8Y7_W2BEG;
	wire [7:0] Tile_X8Y7_W2BEGb;
	wire [15:0] Tile_X8Y7_WW4BEG;
	wire [11:0] Tile_X8Y7_W6BEG;
	wire [3:0] Tile_X9Y7_N1BEG;
	wire [7:0] Tile_X9Y7_N2BEG;
	wire [7:0] Tile_X9Y7_N2BEGb;
	wire [15:0] Tile_X9Y7_N4BEG;
	wire [15:0] Tile_X9Y7_NN4BEG;
	wire [3:0] Tile_X9Y7_E1BEG;
	wire [7:0] Tile_X9Y7_E2BEG;
	wire [7:0] Tile_X9Y7_E2BEGb;
	wire [15:0] Tile_X9Y7_EE4BEG;
	wire [11:0] Tile_X9Y7_E6BEG;
	wire [3:0] Tile_X9Y7_S1BEG;
	wire [7:0] Tile_X9Y7_S2BEG;
	wire [7:0] Tile_X9Y7_S2BEGb;
	wire [15:0] Tile_X9Y7_S4BEG;
	wire [15:0] Tile_X9Y7_SS4BEG;
	wire [17:0] Tile_X9Y7_top2bot;
	wire [3:0] Tile_X9Y7_W1BEG;
	wire [7:0] Tile_X9Y7_W2BEG;
	wire [7:0] Tile_X9Y7_W2BEGb;
	wire [15:0] Tile_X9Y7_WW4BEG;
	wire [11:0] Tile_X9Y7_W6BEG;
	wire [3:0] Tile_X10Y7_N1BEG;
	wire [7:0] Tile_X10Y7_N2BEG;
	wire [7:0] Tile_X10Y7_N2BEGb;
	wire [15:0] Tile_X10Y7_N4BEG;
	wire [15:0] Tile_X10Y7_NN4BEG;
	wire [0:0] Tile_X10Y7_Co;
	wire [3:0] Tile_X10Y7_E1BEG;
	wire [7:0] Tile_X10Y7_E2BEG;
	wire [7:0] Tile_X10Y7_E2BEGb;
	wire [15:0] Tile_X10Y7_EE4BEG;
	wire [11:0] Tile_X10Y7_E6BEG;
	wire [3:0] Tile_X10Y7_S1BEG;
	wire [7:0] Tile_X10Y7_S2BEG;
	wire [7:0] Tile_X10Y7_S2BEGb;
	wire [15:0] Tile_X10Y7_S4BEG;
	wire [15:0] Tile_X10Y7_SS4BEG;
	wire [3:0] Tile_X10Y7_W1BEG;
	wire [7:0] Tile_X10Y7_W2BEG;
	wire [7:0] Tile_X10Y7_W2BEGb;
	wire [15:0] Tile_X10Y7_WW4BEG;
	wire [11:0] Tile_X10Y7_W6BEG;
	wire [3:0] Tile_X11Y7_W1BEG;
	wire [7:0] Tile_X11Y7_W2BEG;
	wire [7:0] Tile_X11Y7_W2BEGb;
	wire [15:0] Tile_X11Y7_WW4BEG;
	wire [11:0] Tile_X11Y7_W6BEG;
	wire [3:0] Tile_X4Y8_E1BEG;
	wire [7:0] Tile_X4Y8_E2BEG;
	wire [7:0] Tile_X4Y8_E2BEGb;
	wire [15:0] Tile_X4Y8_EE4BEG;
	wire [11:0] Tile_X4Y8_E6BEG;
	wire [3:0] Tile_X5Y8_N1BEG;
	wire [7:0] Tile_X5Y8_N2BEG;
	wire [7:0] Tile_X5Y8_N2BEGb;
	wire [15:0] Tile_X5Y8_N4BEG;
	wire [15:0] Tile_X5Y8_NN4BEG;
	wire [9:0] Tile_X5Y8_bot2top;
	wire [3:0] Tile_X5Y8_E1BEG;
	wire [7:0] Tile_X5Y8_E2BEG;
	wire [7:0] Tile_X5Y8_E2BEGb;
	wire [15:0] Tile_X5Y8_EE4BEG;
	wire [11:0] Tile_X5Y8_E6BEG;
	wire [3:0] Tile_X5Y8_S1BEG;
	wire [7:0] Tile_X5Y8_S2BEG;
	wire [7:0] Tile_X5Y8_S2BEGb;
	wire [15:0] Tile_X5Y8_S4BEG;
	wire [15:0] Tile_X5Y8_SS4BEG;
	wire [3:0] Tile_X5Y8_W1BEG;
	wire [7:0] Tile_X5Y8_W2BEG;
	wire [7:0] Tile_X5Y8_W2BEGb;
	wire [15:0] Tile_X5Y8_WW4BEG;
	wire [11:0] Tile_X5Y8_W6BEG;
	wire [3:0] Tile_X6Y8_N1BEG;
	wire [7:0] Tile_X6Y8_N2BEG;
	wire [7:0] Tile_X6Y8_N2BEGb;
	wire [15:0] Tile_X6Y8_N4BEG;
	wire [15:0] Tile_X6Y8_NN4BEG;
	wire [0:0] Tile_X6Y8_Co;
	wire [3:0] Tile_X6Y8_E1BEG;
	wire [7:0] Tile_X6Y8_E2BEG;
	wire [7:0] Tile_X6Y8_E2BEGb;
	wire [15:0] Tile_X6Y8_EE4BEG;
	wire [11:0] Tile_X6Y8_E6BEG;
	wire [3:0] Tile_X6Y8_S1BEG;
	wire [7:0] Tile_X6Y8_S2BEG;
	wire [7:0] Tile_X6Y8_S2BEGb;
	wire [15:0] Tile_X6Y8_S4BEG;
	wire [15:0] Tile_X6Y8_SS4BEG;
	wire [3:0] Tile_X6Y8_W1BEG;
	wire [7:0] Tile_X6Y8_W2BEG;
	wire [7:0] Tile_X6Y8_W2BEGb;
	wire [15:0] Tile_X6Y8_WW4BEG;
	wire [11:0] Tile_X6Y8_W6BEG;
	wire [3:0] Tile_X7Y8_N1BEG;
	wire [7:0] Tile_X7Y8_N2BEG;
	wire [7:0] Tile_X7Y8_N2BEGb;
	wire [15:0] Tile_X7Y8_N4BEG;
	wire [15:0] Tile_X7Y8_NN4BEG;
	wire [0:0] Tile_X7Y8_Co;
	wire [3:0] Tile_X7Y8_E1BEG;
	wire [7:0] Tile_X7Y8_E2BEG;
	wire [7:0] Tile_X7Y8_E2BEGb;
	wire [15:0] Tile_X7Y8_EE4BEG;
	wire [11:0] Tile_X7Y8_E6BEG;
	wire [3:0] Tile_X7Y8_S1BEG;
	wire [7:0] Tile_X7Y8_S2BEG;
	wire [7:0] Tile_X7Y8_S2BEGb;
	wire [15:0] Tile_X7Y8_S4BEG;
	wire [15:0] Tile_X7Y8_SS4BEG;
	wire [3:0] Tile_X7Y8_W1BEG;
	wire [7:0] Tile_X7Y8_W2BEG;
	wire [7:0] Tile_X7Y8_W2BEGb;
	wire [15:0] Tile_X7Y8_WW4BEG;
	wire [11:0] Tile_X7Y8_W6BEG;
	wire [3:0] Tile_X8Y8_N1BEG;
	wire [7:0] Tile_X8Y8_N2BEG;
	wire [7:0] Tile_X8Y8_N2BEGb;
	wire [15:0] Tile_X8Y8_N4BEG;
	wire [15:0] Tile_X8Y8_NN4BEG;
	wire [0:0] Tile_X8Y8_Co;
	wire [3:0] Tile_X8Y8_E1BEG;
	wire [7:0] Tile_X8Y8_E2BEG;
	wire [7:0] Tile_X8Y8_E2BEGb;
	wire [15:0] Tile_X8Y8_EE4BEG;
	wire [11:0] Tile_X8Y8_E6BEG;
	wire [3:0] Tile_X8Y8_S1BEG;
	wire [7:0] Tile_X8Y8_S2BEG;
	wire [7:0] Tile_X8Y8_S2BEGb;
	wire [15:0] Tile_X8Y8_S4BEG;
	wire [15:0] Tile_X8Y8_SS4BEG;
	wire [3:0] Tile_X8Y8_W1BEG;
	wire [7:0] Tile_X8Y8_W2BEG;
	wire [7:0] Tile_X8Y8_W2BEGb;
	wire [15:0] Tile_X8Y8_WW4BEG;
	wire [11:0] Tile_X8Y8_W6BEG;
	wire [3:0] Tile_X9Y8_N1BEG;
	wire [7:0] Tile_X9Y8_N2BEG;
	wire [7:0] Tile_X9Y8_N2BEGb;
	wire [15:0] Tile_X9Y8_N4BEG;
	wire [15:0] Tile_X9Y8_NN4BEG;
	wire [9:0] Tile_X9Y8_bot2top;
	wire [3:0] Tile_X9Y8_E1BEG;
	wire [7:0] Tile_X9Y8_E2BEG;
	wire [7:0] Tile_X9Y8_E2BEGb;
	wire [15:0] Tile_X9Y8_EE4BEG;
	wire [11:0] Tile_X9Y8_E6BEG;
	wire [3:0] Tile_X9Y8_S1BEG;
	wire [7:0] Tile_X9Y8_S2BEG;
	wire [7:0] Tile_X9Y8_S2BEGb;
	wire [15:0] Tile_X9Y8_S4BEG;
	wire [15:0] Tile_X9Y8_SS4BEG;
	wire [3:0] Tile_X9Y8_W1BEG;
	wire [7:0] Tile_X9Y8_W2BEG;
	wire [7:0] Tile_X9Y8_W2BEGb;
	wire [15:0] Tile_X9Y8_WW4BEG;
	wire [11:0] Tile_X9Y8_W6BEG;
	wire [3:0] Tile_X10Y8_N1BEG;
	wire [7:0] Tile_X10Y8_N2BEG;
	wire [7:0] Tile_X10Y8_N2BEGb;
	wire [15:0] Tile_X10Y8_N4BEG;
	wire [15:0] Tile_X10Y8_NN4BEG;
	wire [0:0] Tile_X10Y8_Co;
	wire [3:0] Tile_X10Y8_E1BEG;
	wire [7:0] Tile_X10Y8_E2BEG;
	wire [7:0] Tile_X10Y8_E2BEGb;
	wire [15:0] Tile_X10Y8_EE4BEG;
	wire [11:0] Tile_X10Y8_E6BEG;
	wire [3:0] Tile_X10Y8_S1BEG;
	wire [7:0] Tile_X10Y8_S2BEG;
	wire [7:0] Tile_X10Y8_S2BEGb;
	wire [15:0] Tile_X10Y8_S4BEG;
	wire [15:0] Tile_X10Y8_SS4BEG;
	wire [3:0] Tile_X10Y8_W1BEG;
	wire [7:0] Tile_X10Y8_W2BEG;
	wire [7:0] Tile_X10Y8_W2BEGb;
	wire [15:0] Tile_X10Y8_WW4BEG;
	wire [11:0] Tile_X10Y8_W6BEG;
	wire [3:0] Tile_X11Y8_W1BEG;
	wire [7:0] Tile_X11Y8_W2BEG;
	wire [7:0] Tile_X11Y8_W2BEGb;
	wire [15:0] Tile_X11Y8_WW4BEG;
	wire [11:0] Tile_X11Y8_W6BEG;
	wire [3:0] Tile_X1Y9_S1BEG;
	wire [7:0] Tile_X1Y9_S2BEG;
	wire [7:0] Tile_X1Y9_S2BEGb;
	wire [15:0] Tile_X1Y9_S4BEG;
	wire [15:0] Tile_X1Y9_SS4BEG;
	wire [3:0] Tile_X2Y9_S1BEG;
	wire [7:0] Tile_X2Y9_S2BEG;
	wire [7:0] Tile_X2Y9_S2BEGb;
	wire [15:0] Tile_X2Y9_S4BEG;
	wire [15:0] Tile_X2Y9_SS4BEG;
	wire [3:0] Tile_X3Y9_S1BEG;
	wire [7:0] Tile_X3Y9_S2BEG;
	wire [7:0] Tile_X3Y9_S2BEGb;
	wire [15:0] Tile_X3Y9_S4BEG;
	wire [15:0] Tile_X3Y9_SS4BEG;
	wire [3:0] Tile_X4Y9_E1BEG;
	wire [7:0] Tile_X4Y9_E2BEG;
	wire [7:0] Tile_X4Y9_E2BEGb;
	wire [15:0] Tile_X4Y9_EE4BEG;
	wire [11:0] Tile_X4Y9_E6BEG;
	wire [3:0] Tile_X4Y9_S1BEG;
	wire [7:0] Tile_X4Y9_S2BEG;
	wire [7:0] Tile_X4Y9_S2BEGb;
	wire [15:0] Tile_X4Y9_S4BEG;
	wire [15:0] Tile_X4Y9_SS4BEG;
	wire [3:0] Tile_X5Y9_N1BEG;
	wire [7:0] Tile_X5Y9_N2BEG;
	wire [7:0] Tile_X5Y9_N2BEGb;
	wire [15:0] Tile_X5Y9_N4BEG;
	wire [15:0] Tile_X5Y9_NN4BEG;
	wire [3:0] Tile_X5Y9_E1BEG;
	wire [7:0] Tile_X5Y9_E2BEG;
	wire [7:0] Tile_X5Y9_E2BEGb;
	wire [15:0] Tile_X5Y9_EE4BEG;
	wire [11:0] Tile_X5Y9_E6BEG;
	wire [3:0] Tile_X5Y9_S1BEG;
	wire [7:0] Tile_X5Y9_S2BEG;
	wire [7:0] Tile_X5Y9_S2BEGb;
	wire [15:0] Tile_X5Y9_S4BEG;
	wire [15:0] Tile_X5Y9_SS4BEG;
	wire [17:0] Tile_X5Y9_top2bot;
	wire [3:0] Tile_X5Y9_W1BEG;
	wire [7:0] Tile_X5Y9_W2BEG;
	wire [7:0] Tile_X5Y9_W2BEGb;
	wire [15:0] Tile_X5Y9_WW4BEG;
	wire [11:0] Tile_X5Y9_W6BEG;
	wire [3:0] Tile_X6Y9_N1BEG;
	wire [7:0] Tile_X6Y9_N2BEG;
	wire [7:0] Tile_X6Y9_N2BEGb;
	wire [15:0] Tile_X6Y9_N4BEG;
	wire [15:0] Tile_X6Y9_NN4BEG;
	wire [0:0] Tile_X6Y9_Co;
	wire [3:0] Tile_X6Y9_E1BEG;
	wire [7:0] Tile_X6Y9_E2BEG;
	wire [7:0] Tile_X6Y9_E2BEGb;
	wire [15:0] Tile_X6Y9_EE4BEG;
	wire [11:0] Tile_X6Y9_E6BEG;
	wire [3:0] Tile_X6Y9_S1BEG;
	wire [7:0] Tile_X6Y9_S2BEG;
	wire [7:0] Tile_X6Y9_S2BEGb;
	wire [15:0] Tile_X6Y9_S4BEG;
	wire [15:0] Tile_X6Y9_SS4BEG;
	wire [3:0] Tile_X6Y9_W1BEG;
	wire [7:0] Tile_X6Y9_W2BEG;
	wire [7:0] Tile_X6Y9_W2BEGb;
	wire [15:0] Tile_X6Y9_WW4BEG;
	wire [11:0] Tile_X6Y9_W6BEG;
	wire [3:0] Tile_X7Y9_N1BEG;
	wire [7:0] Tile_X7Y9_N2BEG;
	wire [7:0] Tile_X7Y9_N2BEGb;
	wire [15:0] Tile_X7Y9_N4BEG;
	wire [15:0] Tile_X7Y9_NN4BEG;
	wire [0:0] Tile_X7Y9_Co;
	wire [3:0] Tile_X7Y9_E1BEG;
	wire [7:0] Tile_X7Y9_E2BEG;
	wire [7:0] Tile_X7Y9_E2BEGb;
	wire [15:0] Tile_X7Y9_EE4BEG;
	wire [11:0] Tile_X7Y9_E6BEG;
	wire [3:0] Tile_X7Y9_S1BEG;
	wire [7:0] Tile_X7Y9_S2BEG;
	wire [7:0] Tile_X7Y9_S2BEGb;
	wire [15:0] Tile_X7Y9_S4BEG;
	wire [15:0] Tile_X7Y9_SS4BEG;
	wire [3:0] Tile_X7Y9_W1BEG;
	wire [7:0] Tile_X7Y9_W2BEG;
	wire [7:0] Tile_X7Y9_W2BEGb;
	wire [15:0] Tile_X7Y9_WW4BEG;
	wire [11:0] Tile_X7Y9_W6BEG;
	wire [3:0] Tile_X8Y9_N1BEG;
	wire [7:0] Tile_X8Y9_N2BEG;
	wire [7:0] Tile_X8Y9_N2BEGb;
	wire [15:0] Tile_X8Y9_N4BEG;
	wire [15:0] Tile_X8Y9_NN4BEG;
	wire [0:0] Tile_X8Y9_Co;
	wire [3:0] Tile_X8Y9_E1BEG;
	wire [7:0] Tile_X8Y9_E2BEG;
	wire [7:0] Tile_X8Y9_E2BEGb;
	wire [15:0] Tile_X8Y9_EE4BEG;
	wire [11:0] Tile_X8Y9_E6BEG;
	wire [3:0] Tile_X8Y9_S1BEG;
	wire [7:0] Tile_X8Y9_S2BEG;
	wire [7:0] Tile_X8Y9_S2BEGb;
	wire [15:0] Tile_X8Y9_S4BEG;
	wire [15:0] Tile_X8Y9_SS4BEG;
	wire [3:0] Tile_X8Y9_W1BEG;
	wire [7:0] Tile_X8Y9_W2BEG;
	wire [7:0] Tile_X8Y9_W2BEGb;
	wire [15:0] Tile_X8Y9_WW4BEG;
	wire [11:0] Tile_X8Y9_W6BEG;
	wire [3:0] Tile_X9Y9_N1BEG;
	wire [7:0] Tile_X9Y9_N2BEG;
	wire [7:0] Tile_X9Y9_N2BEGb;
	wire [15:0] Tile_X9Y9_N4BEG;
	wire [15:0] Tile_X9Y9_NN4BEG;
	wire [3:0] Tile_X9Y9_E1BEG;
	wire [7:0] Tile_X9Y9_E2BEG;
	wire [7:0] Tile_X9Y9_E2BEGb;
	wire [15:0] Tile_X9Y9_EE4BEG;
	wire [11:0] Tile_X9Y9_E6BEG;
	wire [3:0] Tile_X9Y9_S1BEG;
	wire [7:0] Tile_X9Y9_S2BEG;
	wire [7:0] Tile_X9Y9_S2BEGb;
	wire [15:0] Tile_X9Y9_S4BEG;
	wire [15:0] Tile_X9Y9_SS4BEG;
	wire [17:0] Tile_X9Y9_top2bot;
	wire [3:0] Tile_X9Y9_W1BEG;
	wire [7:0] Tile_X9Y9_W2BEG;
	wire [7:0] Tile_X9Y9_W2BEGb;
	wire [15:0] Tile_X9Y9_WW4BEG;
	wire [11:0] Tile_X9Y9_W6BEG;
	wire [3:0] Tile_X10Y9_N1BEG;
	wire [7:0] Tile_X10Y9_N2BEG;
	wire [7:0] Tile_X10Y9_N2BEGb;
	wire [15:0] Tile_X10Y9_N4BEG;
	wire [15:0] Tile_X10Y9_NN4BEG;
	wire [0:0] Tile_X10Y9_Co;
	wire [3:0] Tile_X10Y9_E1BEG;
	wire [7:0] Tile_X10Y9_E2BEG;
	wire [7:0] Tile_X10Y9_E2BEGb;
	wire [15:0] Tile_X10Y9_EE4BEG;
	wire [11:0] Tile_X10Y9_E6BEG;
	wire [3:0] Tile_X10Y9_S1BEG;
	wire [7:0] Tile_X10Y9_S2BEG;
	wire [7:0] Tile_X10Y9_S2BEGb;
	wire [15:0] Tile_X10Y9_S4BEG;
	wire [15:0] Tile_X10Y9_SS4BEG;
	wire [3:0] Tile_X10Y9_W1BEG;
	wire [7:0] Tile_X10Y9_W2BEG;
	wire [7:0] Tile_X10Y9_W2BEGb;
	wire [15:0] Tile_X10Y9_WW4BEG;
	wire [11:0] Tile_X10Y9_W6BEG;
	wire [3:0] Tile_X11Y9_S1BEG;
	wire [7:0] Tile_X11Y9_S2BEG;
	wire [7:0] Tile_X11Y9_S2BEGb;
	wire [15:0] Tile_X11Y9_S4BEG;
	wire [15:0] Tile_X11Y9_SS4BEG;
	wire [3:0] Tile_X11Y9_W1BEG;
	wire [7:0] Tile_X11Y9_W2BEG;
	wire [7:0] Tile_X11Y9_W2BEGb;
	wire [15:0] Tile_X11Y9_WW4BEG;
	wire [11:0] Tile_X11Y9_W6BEG;
	wire [3:0] Tile_X12Y9_S1BEG;
	wire [7:0] Tile_X12Y9_S2BEG;
	wire [7:0] Tile_X12Y9_S2BEGb;
	wire [15:0] Tile_X12Y9_S4BEG;
	wire [15:0] Tile_X12Y9_SS4BEG;
	wire [3:0] Tile_X13Y9_S1BEG;
	wire [7:0] Tile_X13Y9_S2BEG;
	wire [7:0] Tile_X13Y9_S2BEGb;
	wire [15:0] Tile_X13Y9_S4BEG;
	wire [15:0] Tile_X13Y9_SS4BEG;
	wire [3:0] Tile_X14Y9_S1BEG;
	wire [7:0] Tile_X14Y9_S2BEG;
	wire [7:0] Tile_X14Y9_S2BEGb;
	wire [15:0] Tile_X14Y9_S4BEG;
	wire [15:0] Tile_X14Y9_SS4BEG;
	wire [3:0] Tile_X15Y9_S1BEG;
	wire [7:0] Tile_X15Y9_S2BEG;
	wire [7:0] Tile_X15Y9_S2BEGb;
	wire [15:0] Tile_X15Y9_S4BEG;
	wire [3:0] Tile_X0Y10_E1BEG;
	wire [7:0] Tile_X0Y10_E2BEG;
	wire [7:0] Tile_X0Y10_E2BEGb;
	wire [15:0] Tile_X0Y10_EE4BEG;
	wire [11:0] Tile_X0Y10_E6BEG;
	wire [3:0] Tile_X1Y10_N1BEG;
	wire [7:0] Tile_X1Y10_N2BEG;
	wire [7:0] Tile_X1Y10_N2BEGb;
	wire [15:0] Tile_X1Y10_N4BEG;
	wire [15:0] Tile_X1Y10_NN4BEG;
	wire [0:0] Tile_X1Y10_Co;
	wire [3:0] Tile_X1Y10_E1BEG;
	wire [7:0] Tile_X1Y10_E2BEG;
	wire [7:0] Tile_X1Y10_E2BEGb;
	wire [15:0] Tile_X1Y10_EE4BEG;
	wire [11:0] Tile_X1Y10_E6BEG;
	wire [3:0] Tile_X1Y10_S1BEG;
	wire [7:0] Tile_X1Y10_S2BEG;
	wire [7:0] Tile_X1Y10_S2BEGb;
	wire [15:0] Tile_X1Y10_S4BEG;
	wire [15:0] Tile_X1Y10_SS4BEG;
	wire [3:0] Tile_X1Y10_W1BEG;
	wire [7:0] Tile_X1Y10_W2BEG;
	wire [7:0] Tile_X1Y10_W2BEGb;
	wire [15:0] Tile_X1Y10_WW4BEG;
	wire [11:0] Tile_X1Y10_W6BEG;
	wire [3:0] Tile_X2Y10_N1BEG;
	wire [7:0] Tile_X2Y10_N2BEG;
	wire [7:0] Tile_X2Y10_N2BEGb;
	wire [15:0] Tile_X2Y10_N4BEG;
	wire [15:0] Tile_X2Y10_NN4BEG;
	wire [3:0] Tile_X2Y10_E1BEG;
	wire [7:0] Tile_X2Y10_E2BEG;
	wire [7:0] Tile_X2Y10_E2BEGb;
	wire [15:0] Tile_X2Y10_EE4BEG;
	wire [11:0] Tile_X2Y10_E6BEG;
	wire [3:0] Tile_X2Y10_S1BEG;
	wire [7:0] Tile_X2Y10_S2BEG;
	wire [7:0] Tile_X2Y10_S2BEGb;
	wire [15:0] Tile_X2Y10_S4BEG;
	wire [15:0] Tile_X2Y10_SS4BEG;
	wire [3:0] Tile_X2Y10_W1BEG;
	wire [7:0] Tile_X2Y10_W2BEG;
	wire [7:0] Tile_X2Y10_W2BEGb;
	wire [15:0] Tile_X2Y10_WW4BEG;
	wire [11:0] Tile_X2Y10_W6BEG;
	wire [3:0] Tile_X3Y10_N1BEG;
	wire [7:0] Tile_X3Y10_N2BEG;
	wire [7:0] Tile_X3Y10_N2BEGb;
	wire [15:0] Tile_X3Y10_N4BEG;
	wire [15:0] Tile_X3Y10_NN4BEG;
	wire [0:0] Tile_X3Y10_Co;
	wire [3:0] Tile_X3Y10_E1BEG;
	wire [7:0] Tile_X3Y10_E2BEG;
	wire [7:0] Tile_X3Y10_E2BEGb;
	wire [15:0] Tile_X3Y10_EE4BEG;
	wire [11:0] Tile_X3Y10_E6BEG;
	wire [3:0] Tile_X3Y10_S1BEG;
	wire [7:0] Tile_X3Y10_S2BEG;
	wire [7:0] Tile_X3Y10_S2BEGb;
	wire [15:0] Tile_X3Y10_S4BEG;
	wire [15:0] Tile_X3Y10_SS4BEG;
	wire [3:0] Tile_X3Y10_W1BEG;
	wire [7:0] Tile_X3Y10_W2BEG;
	wire [7:0] Tile_X3Y10_W2BEGb;
	wire [15:0] Tile_X3Y10_WW4BEG;
	wire [11:0] Tile_X3Y10_W6BEG;
	wire [3:0] Tile_X4Y10_N1BEG;
	wire [7:0] Tile_X4Y10_N2BEG;
	wire [7:0] Tile_X4Y10_N2BEGb;
	wire [15:0] Tile_X4Y10_N4BEG;
	wire [15:0] Tile_X4Y10_NN4BEG;
	wire [0:0] Tile_X4Y10_Co;
	wire [3:0] Tile_X4Y10_E1BEG;
	wire [7:0] Tile_X4Y10_E2BEG;
	wire [7:0] Tile_X4Y10_E2BEGb;
	wire [15:0] Tile_X4Y10_EE4BEG;
	wire [11:0] Tile_X4Y10_E6BEG;
	wire [3:0] Tile_X4Y10_S1BEG;
	wire [7:0] Tile_X4Y10_S2BEG;
	wire [7:0] Tile_X4Y10_S2BEGb;
	wire [15:0] Tile_X4Y10_S4BEG;
	wire [15:0] Tile_X4Y10_SS4BEG;
	wire [3:0] Tile_X4Y10_W1BEG;
	wire [7:0] Tile_X4Y10_W2BEG;
	wire [7:0] Tile_X4Y10_W2BEGb;
	wire [15:0] Tile_X4Y10_WW4BEG;
	wire [11:0] Tile_X4Y10_W6BEG;
	wire [3:0] Tile_X5Y10_N1BEG;
	wire [7:0] Tile_X5Y10_N2BEG;
	wire [7:0] Tile_X5Y10_N2BEGb;
	wire [15:0] Tile_X5Y10_N4BEG;
	wire [15:0] Tile_X5Y10_NN4BEG;
	wire [9:0] Tile_X5Y10_bot2top;
	wire [3:0] Tile_X5Y10_E1BEG;
	wire [7:0] Tile_X5Y10_E2BEG;
	wire [7:0] Tile_X5Y10_E2BEGb;
	wire [15:0] Tile_X5Y10_EE4BEG;
	wire [11:0] Tile_X5Y10_E6BEG;
	wire [3:0] Tile_X5Y10_S1BEG;
	wire [7:0] Tile_X5Y10_S2BEG;
	wire [7:0] Tile_X5Y10_S2BEGb;
	wire [15:0] Tile_X5Y10_S4BEG;
	wire [15:0] Tile_X5Y10_SS4BEG;
	wire [3:0] Tile_X5Y10_W1BEG;
	wire [7:0] Tile_X5Y10_W2BEG;
	wire [7:0] Tile_X5Y10_W2BEGb;
	wire [15:0] Tile_X5Y10_WW4BEG;
	wire [11:0] Tile_X5Y10_W6BEG;
	wire [3:0] Tile_X6Y10_N1BEG;
	wire [7:0] Tile_X6Y10_N2BEG;
	wire [7:0] Tile_X6Y10_N2BEGb;
	wire [15:0] Tile_X6Y10_N4BEG;
	wire [15:0] Tile_X6Y10_NN4BEG;
	wire [0:0] Tile_X6Y10_Co;
	wire [3:0] Tile_X6Y10_E1BEG;
	wire [7:0] Tile_X6Y10_E2BEG;
	wire [7:0] Tile_X6Y10_E2BEGb;
	wire [15:0] Tile_X6Y10_EE4BEG;
	wire [11:0] Tile_X6Y10_E6BEG;
	wire [3:0] Tile_X6Y10_S1BEG;
	wire [7:0] Tile_X6Y10_S2BEG;
	wire [7:0] Tile_X6Y10_S2BEGb;
	wire [15:0] Tile_X6Y10_S4BEG;
	wire [15:0] Tile_X6Y10_SS4BEG;
	wire [3:0] Tile_X6Y10_W1BEG;
	wire [7:0] Tile_X6Y10_W2BEG;
	wire [7:0] Tile_X6Y10_W2BEGb;
	wire [15:0] Tile_X6Y10_WW4BEG;
	wire [11:0] Tile_X6Y10_W6BEG;
	wire [3:0] Tile_X7Y10_N1BEG;
	wire [7:0] Tile_X7Y10_N2BEG;
	wire [7:0] Tile_X7Y10_N2BEGb;
	wire [15:0] Tile_X7Y10_N4BEG;
	wire [15:0] Tile_X7Y10_NN4BEG;
	wire [0:0] Tile_X7Y10_Co;
	wire [3:0] Tile_X7Y10_E1BEG;
	wire [7:0] Tile_X7Y10_E2BEG;
	wire [7:0] Tile_X7Y10_E2BEGb;
	wire [15:0] Tile_X7Y10_EE4BEG;
	wire [11:0] Tile_X7Y10_E6BEG;
	wire [3:0] Tile_X7Y10_S1BEG;
	wire [7:0] Tile_X7Y10_S2BEG;
	wire [7:0] Tile_X7Y10_S2BEGb;
	wire [15:0] Tile_X7Y10_S4BEG;
	wire [15:0] Tile_X7Y10_SS4BEG;
	wire [3:0] Tile_X7Y10_W1BEG;
	wire [7:0] Tile_X7Y10_W2BEG;
	wire [7:0] Tile_X7Y10_W2BEGb;
	wire [15:0] Tile_X7Y10_WW4BEG;
	wire [11:0] Tile_X7Y10_W6BEG;
	wire [3:0] Tile_X8Y10_N1BEG;
	wire [7:0] Tile_X8Y10_N2BEG;
	wire [7:0] Tile_X8Y10_N2BEGb;
	wire [15:0] Tile_X8Y10_N4BEG;
	wire [15:0] Tile_X8Y10_NN4BEG;
	wire [0:0] Tile_X8Y10_Co;
	wire [3:0] Tile_X8Y10_E1BEG;
	wire [7:0] Tile_X8Y10_E2BEG;
	wire [7:0] Tile_X8Y10_E2BEGb;
	wire [15:0] Tile_X8Y10_EE4BEG;
	wire [11:0] Tile_X8Y10_E6BEG;
	wire [3:0] Tile_X8Y10_S1BEG;
	wire [7:0] Tile_X8Y10_S2BEG;
	wire [7:0] Tile_X8Y10_S2BEGb;
	wire [15:0] Tile_X8Y10_S4BEG;
	wire [15:0] Tile_X8Y10_SS4BEG;
	wire [3:0] Tile_X8Y10_W1BEG;
	wire [7:0] Tile_X8Y10_W2BEG;
	wire [7:0] Tile_X8Y10_W2BEGb;
	wire [15:0] Tile_X8Y10_WW4BEG;
	wire [11:0] Tile_X8Y10_W6BEG;
	wire [3:0] Tile_X9Y10_N1BEG;
	wire [7:0] Tile_X9Y10_N2BEG;
	wire [7:0] Tile_X9Y10_N2BEGb;
	wire [15:0] Tile_X9Y10_N4BEG;
	wire [15:0] Tile_X9Y10_NN4BEG;
	wire [9:0] Tile_X9Y10_bot2top;
	wire [3:0] Tile_X9Y10_E1BEG;
	wire [7:0] Tile_X9Y10_E2BEG;
	wire [7:0] Tile_X9Y10_E2BEGb;
	wire [15:0] Tile_X9Y10_EE4BEG;
	wire [11:0] Tile_X9Y10_E6BEG;
	wire [3:0] Tile_X9Y10_S1BEG;
	wire [7:0] Tile_X9Y10_S2BEG;
	wire [7:0] Tile_X9Y10_S2BEGb;
	wire [15:0] Tile_X9Y10_S4BEG;
	wire [15:0] Tile_X9Y10_SS4BEG;
	wire [3:0] Tile_X9Y10_W1BEG;
	wire [7:0] Tile_X9Y10_W2BEG;
	wire [7:0] Tile_X9Y10_W2BEGb;
	wire [15:0] Tile_X9Y10_WW4BEG;
	wire [11:0] Tile_X9Y10_W6BEG;
	wire [3:0] Tile_X10Y10_N1BEG;
	wire [7:0] Tile_X10Y10_N2BEG;
	wire [7:0] Tile_X10Y10_N2BEGb;
	wire [15:0] Tile_X10Y10_N4BEG;
	wire [15:0] Tile_X10Y10_NN4BEG;
	wire [0:0] Tile_X10Y10_Co;
	wire [3:0] Tile_X10Y10_E1BEG;
	wire [7:0] Tile_X10Y10_E2BEG;
	wire [7:0] Tile_X10Y10_E2BEGb;
	wire [15:0] Tile_X10Y10_EE4BEG;
	wire [11:0] Tile_X10Y10_E6BEG;
	wire [3:0] Tile_X10Y10_S1BEG;
	wire [7:0] Tile_X10Y10_S2BEG;
	wire [7:0] Tile_X10Y10_S2BEGb;
	wire [15:0] Tile_X10Y10_S4BEG;
	wire [15:0] Tile_X10Y10_SS4BEG;
	wire [3:0] Tile_X10Y10_W1BEG;
	wire [7:0] Tile_X10Y10_W2BEG;
	wire [7:0] Tile_X10Y10_W2BEGb;
	wire [15:0] Tile_X10Y10_WW4BEG;
	wire [11:0] Tile_X10Y10_W6BEG;
	wire [3:0] Tile_X11Y10_N1BEG;
	wire [7:0] Tile_X11Y10_N2BEG;
	wire [7:0] Tile_X11Y10_N2BEGb;
	wire [15:0] Tile_X11Y10_N4BEG;
	wire [15:0] Tile_X11Y10_NN4BEG;
	wire [0:0] Tile_X11Y10_Co;
	wire [3:0] Tile_X11Y10_E1BEG;
	wire [7:0] Tile_X11Y10_E2BEG;
	wire [7:0] Tile_X11Y10_E2BEGb;
	wire [15:0] Tile_X11Y10_EE4BEG;
	wire [11:0] Tile_X11Y10_E6BEG;
	wire [3:0] Tile_X11Y10_S1BEG;
	wire [7:0] Tile_X11Y10_S2BEG;
	wire [7:0] Tile_X11Y10_S2BEGb;
	wire [15:0] Tile_X11Y10_S4BEG;
	wire [15:0] Tile_X11Y10_SS4BEG;
	wire [3:0] Tile_X11Y10_W1BEG;
	wire [7:0] Tile_X11Y10_W2BEG;
	wire [7:0] Tile_X11Y10_W2BEGb;
	wire [15:0] Tile_X11Y10_WW4BEG;
	wire [11:0] Tile_X11Y10_W6BEG;
	wire [3:0] Tile_X12Y10_N1BEG;
	wire [7:0] Tile_X12Y10_N2BEG;
	wire [7:0] Tile_X12Y10_N2BEGb;
	wire [15:0] Tile_X12Y10_N4BEG;
	wire [15:0] Tile_X12Y10_NN4BEG;
	wire [0:0] Tile_X12Y10_Co;
	wire [3:0] Tile_X12Y10_E1BEG;
	wire [7:0] Tile_X12Y10_E2BEG;
	wire [7:0] Tile_X12Y10_E2BEGb;
	wire [15:0] Tile_X12Y10_EE4BEG;
	wire [11:0] Tile_X12Y10_E6BEG;
	wire [3:0] Tile_X12Y10_S1BEG;
	wire [7:0] Tile_X12Y10_S2BEG;
	wire [7:0] Tile_X12Y10_S2BEGb;
	wire [15:0] Tile_X12Y10_S4BEG;
	wire [15:0] Tile_X12Y10_SS4BEG;
	wire [3:0] Tile_X12Y10_W1BEG;
	wire [7:0] Tile_X12Y10_W2BEG;
	wire [7:0] Tile_X12Y10_W2BEGb;
	wire [15:0] Tile_X12Y10_WW4BEG;
	wire [11:0] Tile_X12Y10_W6BEG;
	wire [3:0] Tile_X13Y10_N1BEG;
	wire [7:0] Tile_X13Y10_N2BEG;
	wire [7:0] Tile_X13Y10_N2BEGb;
	wire [15:0] Tile_X13Y10_N4BEG;
	wire [15:0] Tile_X13Y10_NN4BEG;
	wire [3:0] Tile_X13Y10_E1BEG;
	wire [7:0] Tile_X13Y10_E2BEG;
	wire [7:0] Tile_X13Y10_E2BEGb;
	wire [15:0] Tile_X13Y10_EE4BEG;
	wire [11:0] Tile_X13Y10_E6BEG;
	wire [3:0] Tile_X13Y10_S1BEG;
	wire [7:0] Tile_X13Y10_S2BEG;
	wire [7:0] Tile_X13Y10_S2BEGb;
	wire [15:0] Tile_X13Y10_S4BEG;
	wire [15:0] Tile_X13Y10_SS4BEG;
	wire [3:0] Tile_X13Y10_W1BEG;
	wire [7:0] Tile_X13Y10_W2BEG;
	wire [7:0] Tile_X13Y10_W2BEGb;
	wire [15:0] Tile_X13Y10_WW4BEG;
	wire [11:0] Tile_X13Y10_W6BEG;
	wire [3:0] Tile_X14Y10_N1BEG;
	wire [7:0] Tile_X14Y10_N2BEG;
	wire [7:0] Tile_X14Y10_N2BEGb;
	wire [15:0] Tile_X14Y10_N4BEG;
	wire [15:0] Tile_X14Y10_NN4BEG;
	wire [0:0] Tile_X14Y10_Co;
	wire [3:0] Tile_X14Y10_E1BEG;
	wire [7:0] Tile_X14Y10_E2BEG;
	wire [7:0] Tile_X14Y10_E2BEGb;
	wire [15:0] Tile_X14Y10_EE4BEG;
	wire [11:0] Tile_X14Y10_E6BEG;
	wire [3:0] Tile_X14Y10_S1BEG;
	wire [7:0] Tile_X14Y10_S2BEG;
	wire [7:0] Tile_X14Y10_S2BEGb;
	wire [15:0] Tile_X14Y10_S4BEG;
	wire [15:0] Tile_X14Y10_SS4BEG;
	wire [3:0] Tile_X14Y10_W1BEG;
	wire [7:0] Tile_X14Y10_W2BEG;
	wire [7:0] Tile_X14Y10_W2BEGb;
	wire [15:0] Tile_X14Y10_WW4BEG;
	wire [11:0] Tile_X14Y10_W6BEG;
	wire [3:0] Tile_X15Y10_N1BEG;
	wire [7:0] Tile_X15Y10_N2BEG;
	wire [7:0] Tile_X15Y10_N2BEGb;
	wire [15:0] Tile_X15Y10_N4BEG;
	wire [3:0] Tile_X15Y10_S1BEG;
	wire [7:0] Tile_X15Y10_S2BEG;
	wire [7:0] Tile_X15Y10_S2BEGb;
	wire [15:0] Tile_X15Y10_S4BEG;
	wire [3:0] Tile_X15Y10_W1BEG;
	wire [7:0] Tile_X15Y10_W2BEG;
	wire [7:0] Tile_X15Y10_W2BEGb;
	wire [15:0] Tile_X15Y10_WW4BEG;
	wire [11:0] Tile_X15Y10_W6BEG;
	wire [3:0] Tile_X0Y11_E1BEG;
	wire [7:0] Tile_X0Y11_E2BEG;
	wire [7:0] Tile_X0Y11_E2BEGb;
	wire [15:0] Tile_X0Y11_EE4BEG;
	wire [11:0] Tile_X0Y11_E6BEG;
	wire [3:0] Tile_X1Y11_N1BEG;
	wire [7:0] Tile_X1Y11_N2BEG;
	wire [7:0] Tile_X1Y11_N2BEGb;
	wire [15:0] Tile_X1Y11_N4BEG;
	wire [15:0] Tile_X1Y11_NN4BEG;
	wire [0:0] Tile_X1Y11_Co;
	wire [3:0] Tile_X1Y11_E1BEG;
	wire [7:0] Tile_X1Y11_E2BEG;
	wire [7:0] Tile_X1Y11_E2BEGb;
	wire [15:0] Tile_X1Y11_EE4BEG;
	wire [11:0] Tile_X1Y11_E6BEG;
	wire [3:0] Tile_X1Y11_S1BEG;
	wire [7:0] Tile_X1Y11_S2BEG;
	wire [7:0] Tile_X1Y11_S2BEGb;
	wire [15:0] Tile_X1Y11_S4BEG;
	wire [15:0] Tile_X1Y11_SS4BEG;
	wire [3:0] Tile_X1Y11_W1BEG;
	wire [7:0] Tile_X1Y11_W2BEG;
	wire [7:0] Tile_X1Y11_W2BEGb;
	wire [15:0] Tile_X1Y11_WW4BEG;
	wire [11:0] Tile_X1Y11_W6BEG;
	wire [3:0] Tile_X2Y11_N1BEG;
	wire [7:0] Tile_X2Y11_N2BEG;
	wire [7:0] Tile_X2Y11_N2BEGb;
	wire [15:0] Tile_X2Y11_N4BEG;
	wire [15:0] Tile_X2Y11_NN4BEG;
	wire [3:0] Tile_X2Y11_E1BEG;
	wire [7:0] Tile_X2Y11_E2BEG;
	wire [7:0] Tile_X2Y11_E2BEGb;
	wire [15:0] Tile_X2Y11_EE4BEG;
	wire [11:0] Tile_X2Y11_E6BEG;
	wire [3:0] Tile_X2Y11_S1BEG;
	wire [7:0] Tile_X2Y11_S2BEG;
	wire [7:0] Tile_X2Y11_S2BEGb;
	wire [15:0] Tile_X2Y11_S4BEG;
	wire [15:0] Tile_X2Y11_SS4BEG;
	wire [3:0] Tile_X2Y11_W1BEG;
	wire [7:0] Tile_X2Y11_W2BEG;
	wire [7:0] Tile_X2Y11_W2BEGb;
	wire [15:0] Tile_X2Y11_WW4BEG;
	wire [11:0] Tile_X2Y11_W6BEG;
	wire [3:0] Tile_X3Y11_N1BEG;
	wire [7:0] Tile_X3Y11_N2BEG;
	wire [7:0] Tile_X3Y11_N2BEGb;
	wire [15:0] Tile_X3Y11_N4BEG;
	wire [15:0] Tile_X3Y11_NN4BEG;
	wire [0:0] Tile_X3Y11_Co;
	wire [3:0] Tile_X3Y11_E1BEG;
	wire [7:0] Tile_X3Y11_E2BEG;
	wire [7:0] Tile_X3Y11_E2BEGb;
	wire [15:0] Tile_X3Y11_EE4BEG;
	wire [11:0] Tile_X3Y11_E6BEG;
	wire [3:0] Tile_X3Y11_S1BEG;
	wire [7:0] Tile_X3Y11_S2BEG;
	wire [7:0] Tile_X3Y11_S2BEGb;
	wire [15:0] Tile_X3Y11_S4BEG;
	wire [15:0] Tile_X3Y11_SS4BEG;
	wire [3:0] Tile_X3Y11_W1BEG;
	wire [7:0] Tile_X3Y11_W2BEG;
	wire [7:0] Tile_X3Y11_W2BEGb;
	wire [15:0] Tile_X3Y11_WW4BEG;
	wire [11:0] Tile_X3Y11_W6BEG;
	wire [3:0] Tile_X4Y11_N1BEG;
	wire [7:0] Tile_X4Y11_N2BEG;
	wire [7:0] Tile_X4Y11_N2BEGb;
	wire [15:0] Tile_X4Y11_N4BEG;
	wire [15:0] Tile_X4Y11_NN4BEG;
	wire [0:0] Tile_X4Y11_Co;
	wire [3:0] Tile_X4Y11_E1BEG;
	wire [7:0] Tile_X4Y11_E2BEG;
	wire [7:0] Tile_X4Y11_E2BEGb;
	wire [15:0] Tile_X4Y11_EE4BEG;
	wire [11:0] Tile_X4Y11_E6BEG;
	wire [3:0] Tile_X4Y11_S1BEG;
	wire [7:0] Tile_X4Y11_S2BEG;
	wire [7:0] Tile_X4Y11_S2BEGb;
	wire [15:0] Tile_X4Y11_S4BEG;
	wire [15:0] Tile_X4Y11_SS4BEG;
	wire [3:0] Tile_X4Y11_W1BEG;
	wire [7:0] Tile_X4Y11_W2BEG;
	wire [7:0] Tile_X4Y11_W2BEGb;
	wire [15:0] Tile_X4Y11_WW4BEG;
	wire [11:0] Tile_X4Y11_W6BEG;
	wire [3:0] Tile_X5Y11_N1BEG;
	wire [7:0] Tile_X5Y11_N2BEG;
	wire [7:0] Tile_X5Y11_N2BEGb;
	wire [15:0] Tile_X5Y11_N4BEG;
	wire [15:0] Tile_X5Y11_NN4BEG;
	wire [3:0] Tile_X5Y11_E1BEG;
	wire [7:0] Tile_X5Y11_E2BEG;
	wire [7:0] Tile_X5Y11_E2BEGb;
	wire [15:0] Tile_X5Y11_EE4BEG;
	wire [11:0] Tile_X5Y11_E6BEG;
	wire [3:0] Tile_X5Y11_S1BEG;
	wire [7:0] Tile_X5Y11_S2BEG;
	wire [7:0] Tile_X5Y11_S2BEGb;
	wire [15:0] Tile_X5Y11_S4BEG;
	wire [15:0] Tile_X5Y11_SS4BEG;
	wire [17:0] Tile_X5Y11_top2bot;
	wire [3:0] Tile_X5Y11_W1BEG;
	wire [7:0] Tile_X5Y11_W2BEG;
	wire [7:0] Tile_X5Y11_W2BEGb;
	wire [15:0] Tile_X5Y11_WW4BEG;
	wire [11:0] Tile_X5Y11_W6BEG;
	wire [3:0] Tile_X6Y11_N1BEG;
	wire [7:0] Tile_X6Y11_N2BEG;
	wire [7:0] Tile_X6Y11_N2BEGb;
	wire [15:0] Tile_X6Y11_N4BEG;
	wire [15:0] Tile_X6Y11_NN4BEG;
	wire [0:0] Tile_X6Y11_Co;
	wire [3:0] Tile_X6Y11_E1BEG;
	wire [7:0] Tile_X6Y11_E2BEG;
	wire [7:0] Tile_X6Y11_E2BEGb;
	wire [15:0] Tile_X6Y11_EE4BEG;
	wire [11:0] Tile_X6Y11_E6BEG;
	wire [3:0] Tile_X6Y11_S1BEG;
	wire [7:0] Tile_X6Y11_S2BEG;
	wire [7:0] Tile_X6Y11_S2BEGb;
	wire [15:0] Tile_X6Y11_S4BEG;
	wire [15:0] Tile_X6Y11_SS4BEG;
	wire [3:0] Tile_X6Y11_W1BEG;
	wire [7:0] Tile_X6Y11_W2BEG;
	wire [7:0] Tile_X6Y11_W2BEGb;
	wire [15:0] Tile_X6Y11_WW4BEG;
	wire [11:0] Tile_X6Y11_W6BEG;
	wire [3:0] Tile_X7Y11_N1BEG;
	wire [7:0] Tile_X7Y11_N2BEG;
	wire [7:0] Tile_X7Y11_N2BEGb;
	wire [15:0] Tile_X7Y11_N4BEG;
	wire [15:0] Tile_X7Y11_NN4BEG;
	wire [0:0] Tile_X7Y11_Co;
	wire [3:0] Tile_X7Y11_E1BEG;
	wire [7:0] Tile_X7Y11_E2BEG;
	wire [7:0] Tile_X7Y11_E2BEGb;
	wire [15:0] Tile_X7Y11_EE4BEG;
	wire [11:0] Tile_X7Y11_E6BEG;
	wire [3:0] Tile_X7Y11_S1BEG;
	wire [7:0] Tile_X7Y11_S2BEG;
	wire [7:0] Tile_X7Y11_S2BEGb;
	wire [15:0] Tile_X7Y11_S4BEG;
	wire [15:0] Tile_X7Y11_SS4BEG;
	wire [3:0] Tile_X7Y11_W1BEG;
	wire [7:0] Tile_X7Y11_W2BEG;
	wire [7:0] Tile_X7Y11_W2BEGb;
	wire [15:0] Tile_X7Y11_WW4BEG;
	wire [11:0] Tile_X7Y11_W6BEG;
	wire [3:0] Tile_X8Y11_N1BEG;
	wire [7:0] Tile_X8Y11_N2BEG;
	wire [7:0] Tile_X8Y11_N2BEGb;
	wire [15:0] Tile_X8Y11_N4BEG;
	wire [15:0] Tile_X8Y11_NN4BEG;
	wire [0:0] Tile_X8Y11_Co;
	wire [3:0] Tile_X8Y11_E1BEG;
	wire [7:0] Tile_X8Y11_E2BEG;
	wire [7:0] Tile_X8Y11_E2BEGb;
	wire [15:0] Tile_X8Y11_EE4BEG;
	wire [11:0] Tile_X8Y11_E6BEG;
	wire [3:0] Tile_X8Y11_S1BEG;
	wire [7:0] Tile_X8Y11_S2BEG;
	wire [7:0] Tile_X8Y11_S2BEGb;
	wire [15:0] Tile_X8Y11_S4BEG;
	wire [15:0] Tile_X8Y11_SS4BEG;
	wire [3:0] Tile_X8Y11_W1BEG;
	wire [7:0] Tile_X8Y11_W2BEG;
	wire [7:0] Tile_X8Y11_W2BEGb;
	wire [15:0] Tile_X8Y11_WW4BEG;
	wire [11:0] Tile_X8Y11_W6BEG;
	wire [3:0] Tile_X9Y11_N1BEG;
	wire [7:0] Tile_X9Y11_N2BEG;
	wire [7:0] Tile_X9Y11_N2BEGb;
	wire [15:0] Tile_X9Y11_N4BEG;
	wire [15:0] Tile_X9Y11_NN4BEG;
	wire [3:0] Tile_X9Y11_E1BEG;
	wire [7:0] Tile_X9Y11_E2BEG;
	wire [7:0] Tile_X9Y11_E2BEGb;
	wire [15:0] Tile_X9Y11_EE4BEG;
	wire [11:0] Tile_X9Y11_E6BEG;
	wire [3:0] Tile_X9Y11_S1BEG;
	wire [7:0] Tile_X9Y11_S2BEG;
	wire [7:0] Tile_X9Y11_S2BEGb;
	wire [15:0] Tile_X9Y11_S4BEG;
	wire [15:0] Tile_X9Y11_SS4BEG;
	wire [17:0] Tile_X9Y11_top2bot;
	wire [3:0] Tile_X9Y11_W1BEG;
	wire [7:0] Tile_X9Y11_W2BEG;
	wire [7:0] Tile_X9Y11_W2BEGb;
	wire [15:0] Tile_X9Y11_WW4BEG;
	wire [11:0] Tile_X9Y11_W6BEG;
	wire [3:0] Tile_X10Y11_N1BEG;
	wire [7:0] Tile_X10Y11_N2BEG;
	wire [7:0] Tile_X10Y11_N2BEGb;
	wire [15:0] Tile_X10Y11_N4BEG;
	wire [15:0] Tile_X10Y11_NN4BEG;
	wire [0:0] Tile_X10Y11_Co;
	wire [3:0] Tile_X10Y11_E1BEG;
	wire [7:0] Tile_X10Y11_E2BEG;
	wire [7:0] Tile_X10Y11_E2BEGb;
	wire [15:0] Tile_X10Y11_EE4BEG;
	wire [11:0] Tile_X10Y11_E6BEG;
	wire [3:0] Tile_X10Y11_S1BEG;
	wire [7:0] Tile_X10Y11_S2BEG;
	wire [7:0] Tile_X10Y11_S2BEGb;
	wire [15:0] Tile_X10Y11_S4BEG;
	wire [15:0] Tile_X10Y11_SS4BEG;
	wire [3:0] Tile_X10Y11_W1BEG;
	wire [7:0] Tile_X10Y11_W2BEG;
	wire [7:0] Tile_X10Y11_W2BEGb;
	wire [15:0] Tile_X10Y11_WW4BEG;
	wire [11:0] Tile_X10Y11_W6BEG;
	wire [3:0] Tile_X11Y11_N1BEG;
	wire [7:0] Tile_X11Y11_N2BEG;
	wire [7:0] Tile_X11Y11_N2BEGb;
	wire [15:0] Tile_X11Y11_N4BEG;
	wire [15:0] Tile_X11Y11_NN4BEG;
	wire [0:0] Tile_X11Y11_Co;
	wire [3:0] Tile_X11Y11_E1BEG;
	wire [7:0] Tile_X11Y11_E2BEG;
	wire [7:0] Tile_X11Y11_E2BEGb;
	wire [15:0] Tile_X11Y11_EE4BEG;
	wire [11:0] Tile_X11Y11_E6BEG;
	wire [3:0] Tile_X11Y11_S1BEG;
	wire [7:0] Tile_X11Y11_S2BEG;
	wire [7:0] Tile_X11Y11_S2BEGb;
	wire [15:0] Tile_X11Y11_S4BEG;
	wire [15:0] Tile_X11Y11_SS4BEG;
	wire [3:0] Tile_X11Y11_W1BEG;
	wire [7:0] Tile_X11Y11_W2BEG;
	wire [7:0] Tile_X11Y11_W2BEGb;
	wire [15:0] Tile_X11Y11_WW4BEG;
	wire [11:0] Tile_X11Y11_W6BEG;
	wire [3:0] Tile_X12Y11_N1BEG;
	wire [7:0] Tile_X12Y11_N2BEG;
	wire [7:0] Tile_X12Y11_N2BEGb;
	wire [15:0] Tile_X12Y11_N4BEG;
	wire [15:0] Tile_X12Y11_NN4BEG;
	wire [0:0] Tile_X12Y11_Co;
	wire [3:0] Tile_X12Y11_E1BEG;
	wire [7:0] Tile_X12Y11_E2BEG;
	wire [7:0] Tile_X12Y11_E2BEGb;
	wire [15:0] Tile_X12Y11_EE4BEG;
	wire [11:0] Tile_X12Y11_E6BEG;
	wire [3:0] Tile_X12Y11_S1BEG;
	wire [7:0] Tile_X12Y11_S2BEG;
	wire [7:0] Tile_X12Y11_S2BEGb;
	wire [15:0] Tile_X12Y11_S4BEG;
	wire [15:0] Tile_X12Y11_SS4BEG;
	wire [3:0] Tile_X12Y11_W1BEG;
	wire [7:0] Tile_X12Y11_W2BEG;
	wire [7:0] Tile_X12Y11_W2BEGb;
	wire [15:0] Tile_X12Y11_WW4BEG;
	wire [11:0] Tile_X12Y11_W6BEG;
	wire [3:0] Tile_X13Y11_N1BEG;
	wire [7:0] Tile_X13Y11_N2BEG;
	wire [7:0] Tile_X13Y11_N2BEGb;
	wire [15:0] Tile_X13Y11_N4BEG;
	wire [15:0] Tile_X13Y11_NN4BEG;
	wire [3:0] Tile_X13Y11_E1BEG;
	wire [7:0] Tile_X13Y11_E2BEG;
	wire [7:0] Tile_X13Y11_E2BEGb;
	wire [15:0] Tile_X13Y11_EE4BEG;
	wire [11:0] Tile_X13Y11_E6BEG;
	wire [3:0] Tile_X13Y11_S1BEG;
	wire [7:0] Tile_X13Y11_S2BEG;
	wire [7:0] Tile_X13Y11_S2BEGb;
	wire [15:0] Tile_X13Y11_S4BEG;
	wire [15:0] Tile_X13Y11_SS4BEG;
	wire [3:0] Tile_X13Y11_W1BEG;
	wire [7:0] Tile_X13Y11_W2BEG;
	wire [7:0] Tile_X13Y11_W2BEGb;
	wire [15:0] Tile_X13Y11_WW4BEG;
	wire [11:0] Tile_X13Y11_W6BEG;
	wire [3:0] Tile_X14Y11_N1BEG;
	wire [7:0] Tile_X14Y11_N2BEG;
	wire [7:0] Tile_X14Y11_N2BEGb;
	wire [15:0] Tile_X14Y11_N4BEG;
	wire [15:0] Tile_X14Y11_NN4BEG;
	wire [0:0] Tile_X14Y11_Co;
	wire [3:0] Tile_X14Y11_E1BEG;
	wire [7:0] Tile_X14Y11_E2BEG;
	wire [7:0] Tile_X14Y11_E2BEGb;
	wire [15:0] Tile_X14Y11_EE4BEG;
	wire [11:0] Tile_X14Y11_E6BEG;
	wire [3:0] Tile_X14Y11_S1BEG;
	wire [7:0] Tile_X14Y11_S2BEG;
	wire [7:0] Tile_X14Y11_S2BEGb;
	wire [15:0] Tile_X14Y11_S4BEG;
	wire [15:0] Tile_X14Y11_SS4BEG;
	wire [3:0] Tile_X14Y11_W1BEG;
	wire [7:0] Tile_X14Y11_W2BEG;
	wire [7:0] Tile_X14Y11_W2BEGb;
	wire [15:0] Tile_X14Y11_WW4BEG;
	wire [11:0] Tile_X14Y11_W6BEG;
	wire [3:0] Tile_X15Y11_N1BEG;
	wire [7:0] Tile_X15Y11_N2BEG;
	wire [7:0] Tile_X15Y11_N2BEGb;
	wire [15:0] Tile_X15Y11_N4BEG;
	wire [3:0] Tile_X15Y11_S1BEG;
	wire [7:0] Tile_X15Y11_S2BEG;
	wire [7:0] Tile_X15Y11_S2BEGb;
	wire [15:0] Tile_X15Y11_S4BEG;
	wire [3:0] Tile_X15Y11_W1BEG;
	wire [7:0] Tile_X15Y11_W2BEG;
	wire [7:0] Tile_X15Y11_W2BEGb;
	wire [15:0] Tile_X15Y11_WW4BEG;
	wire [11:0] Tile_X15Y11_W6BEG;
	wire [3:0] Tile_X0Y12_E1BEG;
	wire [7:0] Tile_X0Y12_E2BEG;
	wire [7:0] Tile_X0Y12_E2BEGb;
	wire [15:0] Tile_X0Y12_EE4BEG;
	wire [11:0] Tile_X0Y12_E6BEG;
	wire [3:0] Tile_X1Y12_N1BEG;
	wire [7:0] Tile_X1Y12_N2BEG;
	wire [7:0] Tile_X1Y12_N2BEGb;
	wire [15:0] Tile_X1Y12_N4BEG;
	wire [15:0] Tile_X1Y12_NN4BEG;
	wire [0:0] Tile_X1Y12_Co;
	wire [3:0] Tile_X1Y12_E1BEG;
	wire [7:0] Tile_X1Y12_E2BEG;
	wire [7:0] Tile_X1Y12_E2BEGb;
	wire [15:0] Tile_X1Y12_EE4BEG;
	wire [11:0] Tile_X1Y12_E6BEG;
	wire [3:0] Tile_X1Y12_S1BEG;
	wire [7:0] Tile_X1Y12_S2BEG;
	wire [7:0] Tile_X1Y12_S2BEGb;
	wire [15:0] Tile_X1Y12_S4BEG;
	wire [15:0] Tile_X1Y12_SS4BEG;
	wire [3:0] Tile_X1Y12_W1BEG;
	wire [7:0] Tile_X1Y12_W2BEG;
	wire [7:0] Tile_X1Y12_W2BEGb;
	wire [15:0] Tile_X1Y12_WW4BEG;
	wire [11:0] Tile_X1Y12_W6BEG;
	wire [3:0] Tile_X2Y12_N1BEG;
	wire [7:0] Tile_X2Y12_N2BEG;
	wire [7:0] Tile_X2Y12_N2BEGb;
	wire [15:0] Tile_X2Y12_N4BEG;
	wire [15:0] Tile_X2Y12_NN4BEG;
	wire [3:0] Tile_X2Y12_E1BEG;
	wire [7:0] Tile_X2Y12_E2BEG;
	wire [7:0] Tile_X2Y12_E2BEGb;
	wire [15:0] Tile_X2Y12_EE4BEG;
	wire [11:0] Tile_X2Y12_E6BEG;
	wire [3:0] Tile_X2Y12_S1BEG;
	wire [7:0] Tile_X2Y12_S2BEG;
	wire [7:0] Tile_X2Y12_S2BEGb;
	wire [15:0] Tile_X2Y12_S4BEG;
	wire [15:0] Tile_X2Y12_SS4BEG;
	wire [3:0] Tile_X2Y12_W1BEG;
	wire [7:0] Tile_X2Y12_W2BEG;
	wire [7:0] Tile_X2Y12_W2BEGb;
	wire [15:0] Tile_X2Y12_WW4BEG;
	wire [11:0] Tile_X2Y12_W6BEG;
	wire [3:0] Tile_X3Y12_N1BEG;
	wire [7:0] Tile_X3Y12_N2BEG;
	wire [7:0] Tile_X3Y12_N2BEGb;
	wire [15:0] Tile_X3Y12_N4BEG;
	wire [15:0] Tile_X3Y12_NN4BEG;
	wire [0:0] Tile_X3Y12_Co;
	wire [3:0] Tile_X3Y12_E1BEG;
	wire [7:0] Tile_X3Y12_E2BEG;
	wire [7:0] Tile_X3Y12_E2BEGb;
	wire [15:0] Tile_X3Y12_EE4BEG;
	wire [11:0] Tile_X3Y12_E6BEG;
	wire [3:0] Tile_X3Y12_S1BEG;
	wire [7:0] Tile_X3Y12_S2BEG;
	wire [7:0] Tile_X3Y12_S2BEGb;
	wire [15:0] Tile_X3Y12_S4BEG;
	wire [15:0] Tile_X3Y12_SS4BEG;
	wire [3:0] Tile_X3Y12_W1BEG;
	wire [7:0] Tile_X3Y12_W2BEG;
	wire [7:0] Tile_X3Y12_W2BEGb;
	wire [15:0] Tile_X3Y12_WW4BEG;
	wire [11:0] Tile_X3Y12_W6BEG;
	wire [3:0] Tile_X4Y12_N1BEG;
	wire [7:0] Tile_X4Y12_N2BEG;
	wire [7:0] Tile_X4Y12_N2BEGb;
	wire [15:0] Tile_X4Y12_N4BEG;
	wire [15:0] Tile_X4Y12_NN4BEG;
	wire [0:0] Tile_X4Y12_Co;
	wire [3:0] Tile_X4Y12_E1BEG;
	wire [7:0] Tile_X4Y12_E2BEG;
	wire [7:0] Tile_X4Y12_E2BEGb;
	wire [15:0] Tile_X4Y12_EE4BEG;
	wire [11:0] Tile_X4Y12_E6BEG;
	wire [3:0] Tile_X4Y12_S1BEG;
	wire [7:0] Tile_X4Y12_S2BEG;
	wire [7:0] Tile_X4Y12_S2BEGb;
	wire [15:0] Tile_X4Y12_S4BEG;
	wire [15:0] Tile_X4Y12_SS4BEG;
	wire [3:0] Tile_X4Y12_W1BEG;
	wire [7:0] Tile_X4Y12_W2BEG;
	wire [7:0] Tile_X4Y12_W2BEGb;
	wire [15:0] Tile_X4Y12_WW4BEG;
	wire [11:0] Tile_X4Y12_W6BEG;
	wire [3:0] Tile_X5Y12_N1BEG;
	wire [7:0] Tile_X5Y12_N2BEG;
	wire [7:0] Tile_X5Y12_N2BEGb;
	wire [15:0] Tile_X5Y12_N4BEG;
	wire [15:0] Tile_X5Y12_NN4BEG;
	wire [9:0] Tile_X5Y12_bot2top;
	wire [3:0] Tile_X5Y12_E1BEG;
	wire [7:0] Tile_X5Y12_E2BEG;
	wire [7:0] Tile_X5Y12_E2BEGb;
	wire [15:0] Tile_X5Y12_EE4BEG;
	wire [11:0] Tile_X5Y12_E6BEG;
	wire [3:0] Tile_X5Y12_S1BEG;
	wire [7:0] Tile_X5Y12_S2BEG;
	wire [7:0] Tile_X5Y12_S2BEGb;
	wire [15:0] Tile_X5Y12_S4BEG;
	wire [15:0] Tile_X5Y12_SS4BEG;
	wire [3:0] Tile_X5Y12_W1BEG;
	wire [7:0] Tile_X5Y12_W2BEG;
	wire [7:0] Tile_X5Y12_W2BEGb;
	wire [15:0] Tile_X5Y12_WW4BEG;
	wire [11:0] Tile_X5Y12_W6BEG;
	wire [3:0] Tile_X6Y12_N1BEG;
	wire [7:0] Tile_X6Y12_N2BEG;
	wire [7:0] Tile_X6Y12_N2BEGb;
	wire [15:0] Tile_X6Y12_N4BEG;
	wire [15:0] Tile_X6Y12_NN4BEG;
	wire [0:0] Tile_X6Y12_Co;
	wire [3:0] Tile_X6Y12_E1BEG;
	wire [7:0] Tile_X6Y12_E2BEG;
	wire [7:0] Tile_X6Y12_E2BEGb;
	wire [15:0] Tile_X6Y12_EE4BEG;
	wire [11:0] Tile_X6Y12_E6BEG;
	wire [3:0] Tile_X6Y12_S1BEG;
	wire [7:0] Tile_X6Y12_S2BEG;
	wire [7:0] Tile_X6Y12_S2BEGb;
	wire [15:0] Tile_X6Y12_S4BEG;
	wire [15:0] Tile_X6Y12_SS4BEG;
	wire [3:0] Tile_X6Y12_W1BEG;
	wire [7:0] Tile_X6Y12_W2BEG;
	wire [7:0] Tile_X6Y12_W2BEGb;
	wire [15:0] Tile_X6Y12_WW4BEG;
	wire [11:0] Tile_X6Y12_W6BEG;
	wire [3:0] Tile_X7Y12_N1BEG;
	wire [7:0] Tile_X7Y12_N2BEG;
	wire [7:0] Tile_X7Y12_N2BEGb;
	wire [15:0] Tile_X7Y12_N4BEG;
	wire [15:0] Tile_X7Y12_NN4BEG;
	wire [0:0] Tile_X7Y12_Co;
	wire [3:0] Tile_X7Y12_E1BEG;
	wire [7:0] Tile_X7Y12_E2BEG;
	wire [7:0] Tile_X7Y12_E2BEGb;
	wire [15:0] Tile_X7Y12_EE4BEG;
	wire [11:0] Tile_X7Y12_E6BEG;
	wire [3:0] Tile_X7Y12_S1BEG;
	wire [7:0] Tile_X7Y12_S2BEG;
	wire [7:0] Tile_X7Y12_S2BEGb;
	wire [15:0] Tile_X7Y12_S4BEG;
	wire [15:0] Tile_X7Y12_SS4BEG;
	wire [3:0] Tile_X7Y12_W1BEG;
	wire [7:0] Tile_X7Y12_W2BEG;
	wire [7:0] Tile_X7Y12_W2BEGb;
	wire [15:0] Tile_X7Y12_WW4BEG;
	wire [11:0] Tile_X7Y12_W6BEG;
	wire [3:0] Tile_X8Y12_N1BEG;
	wire [7:0] Tile_X8Y12_N2BEG;
	wire [7:0] Tile_X8Y12_N2BEGb;
	wire [15:0] Tile_X8Y12_N4BEG;
	wire [15:0] Tile_X8Y12_NN4BEG;
	wire [0:0] Tile_X8Y12_Co;
	wire [3:0] Tile_X8Y12_E1BEG;
	wire [7:0] Tile_X8Y12_E2BEG;
	wire [7:0] Tile_X8Y12_E2BEGb;
	wire [15:0] Tile_X8Y12_EE4BEG;
	wire [11:0] Tile_X8Y12_E6BEG;
	wire [3:0] Tile_X8Y12_S1BEG;
	wire [7:0] Tile_X8Y12_S2BEG;
	wire [7:0] Tile_X8Y12_S2BEGb;
	wire [15:0] Tile_X8Y12_S4BEG;
	wire [15:0] Tile_X8Y12_SS4BEG;
	wire [3:0] Tile_X8Y12_W1BEG;
	wire [7:0] Tile_X8Y12_W2BEG;
	wire [7:0] Tile_X8Y12_W2BEGb;
	wire [15:0] Tile_X8Y12_WW4BEG;
	wire [11:0] Tile_X8Y12_W6BEG;
	wire [3:0] Tile_X9Y12_N1BEG;
	wire [7:0] Tile_X9Y12_N2BEG;
	wire [7:0] Tile_X9Y12_N2BEGb;
	wire [15:0] Tile_X9Y12_N4BEG;
	wire [15:0] Tile_X9Y12_NN4BEG;
	wire [9:0] Tile_X9Y12_bot2top;
	wire [3:0] Tile_X9Y12_E1BEG;
	wire [7:0] Tile_X9Y12_E2BEG;
	wire [7:0] Tile_X9Y12_E2BEGb;
	wire [15:0] Tile_X9Y12_EE4BEG;
	wire [11:0] Tile_X9Y12_E6BEG;
	wire [3:0] Tile_X9Y12_S1BEG;
	wire [7:0] Tile_X9Y12_S2BEG;
	wire [7:0] Tile_X9Y12_S2BEGb;
	wire [15:0] Tile_X9Y12_S4BEG;
	wire [15:0] Tile_X9Y12_SS4BEG;
	wire [3:0] Tile_X9Y12_W1BEG;
	wire [7:0] Tile_X9Y12_W2BEG;
	wire [7:0] Tile_X9Y12_W2BEGb;
	wire [15:0] Tile_X9Y12_WW4BEG;
	wire [11:0] Tile_X9Y12_W6BEG;
	wire [3:0] Tile_X10Y12_N1BEG;
	wire [7:0] Tile_X10Y12_N2BEG;
	wire [7:0] Tile_X10Y12_N2BEGb;
	wire [15:0] Tile_X10Y12_N4BEG;
	wire [15:0] Tile_X10Y12_NN4BEG;
	wire [0:0] Tile_X10Y12_Co;
	wire [3:0] Tile_X10Y12_E1BEG;
	wire [7:0] Tile_X10Y12_E2BEG;
	wire [7:0] Tile_X10Y12_E2BEGb;
	wire [15:0] Tile_X10Y12_EE4BEG;
	wire [11:0] Tile_X10Y12_E6BEG;
	wire [3:0] Tile_X10Y12_S1BEG;
	wire [7:0] Tile_X10Y12_S2BEG;
	wire [7:0] Tile_X10Y12_S2BEGb;
	wire [15:0] Tile_X10Y12_S4BEG;
	wire [15:0] Tile_X10Y12_SS4BEG;
	wire [3:0] Tile_X10Y12_W1BEG;
	wire [7:0] Tile_X10Y12_W2BEG;
	wire [7:0] Tile_X10Y12_W2BEGb;
	wire [15:0] Tile_X10Y12_WW4BEG;
	wire [11:0] Tile_X10Y12_W6BEG;
	wire [3:0] Tile_X11Y12_N1BEG;
	wire [7:0] Tile_X11Y12_N2BEG;
	wire [7:0] Tile_X11Y12_N2BEGb;
	wire [15:0] Tile_X11Y12_N4BEG;
	wire [15:0] Tile_X11Y12_NN4BEG;
	wire [0:0] Tile_X11Y12_Co;
	wire [3:0] Tile_X11Y12_E1BEG;
	wire [7:0] Tile_X11Y12_E2BEG;
	wire [7:0] Tile_X11Y12_E2BEGb;
	wire [15:0] Tile_X11Y12_EE4BEG;
	wire [11:0] Tile_X11Y12_E6BEG;
	wire [3:0] Tile_X11Y12_S1BEG;
	wire [7:0] Tile_X11Y12_S2BEG;
	wire [7:0] Tile_X11Y12_S2BEGb;
	wire [15:0] Tile_X11Y12_S4BEG;
	wire [15:0] Tile_X11Y12_SS4BEG;
	wire [3:0] Tile_X11Y12_W1BEG;
	wire [7:0] Tile_X11Y12_W2BEG;
	wire [7:0] Tile_X11Y12_W2BEGb;
	wire [15:0] Tile_X11Y12_WW4BEG;
	wire [11:0] Tile_X11Y12_W6BEG;
	wire [3:0] Tile_X12Y12_N1BEG;
	wire [7:0] Tile_X12Y12_N2BEG;
	wire [7:0] Tile_X12Y12_N2BEGb;
	wire [15:0] Tile_X12Y12_N4BEG;
	wire [15:0] Tile_X12Y12_NN4BEG;
	wire [0:0] Tile_X12Y12_Co;
	wire [3:0] Tile_X12Y12_E1BEG;
	wire [7:0] Tile_X12Y12_E2BEG;
	wire [7:0] Tile_X12Y12_E2BEGb;
	wire [15:0] Tile_X12Y12_EE4BEG;
	wire [11:0] Tile_X12Y12_E6BEG;
	wire [3:0] Tile_X12Y12_S1BEG;
	wire [7:0] Tile_X12Y12_S2BEG;
	wire [7:0] Tile_X12Y12_S2BEGb;
	wire [15:0] Tile_X12Y12_S4BEG;
	wire [15:0] Tile_X12Y12_SS4BEG;
	wire [3:0] Tile_X12Y12_W1BEG;
	wire [7:0] Tile_X12Y12_W2BEG;
	wire [7:0] Tile_X12Y12_W2BEGb;
	wire [15:0] Tile_X12Y12_WW4BEG;
	wire [11:0] Tile_X12Y12_W6BEG;
	wire [3:0] Tile_X13Y12_N1BEG;
	wire [7:0] Tile_X13Y12_N2BEG;
	wire [7:0] Tile_X13Y12_N2BEGb;
	wire [15:0] Tile_X13Y12_N4BEG;
	wire [15:0] Tile_X13Y12_NN4BEG;
	wire [3:0] Tile_X13Y12_E1BEG;
	wire [7:0] Tile_X13Y12_E2BEG;
	wire [7:0] Tile_X13Y12_E2BEGb;
	wire [15:0] Tile_X13Y12_EE4BEG;
	wire [11:0] Tile_X13Y12_E6BEG;
	wire [3:0] Tile_X13Y12_S1BEG;
	wire [7:0] Tile_X13Y12_S2BEG;
	wire [7:0] Tile_X13Y12_S2BEGb;
	wire [15:0] Tile_X13Y12_S4BEG;
	wire [15:0] Tile_X13Y12_SS4BEG;
	wire [3:0] Tile_X13Y12_W1BEG;
	wire [7:0] Tile_X13Y12_W2BEG;
	wire [7:0] Tile_X13Y12_W2BEGb;
	wire [15:0] Tile_X13Y12_WW4BEG;
	wire [11:0] Tile_X13Y12_W6BEG;
	wire [3:0] Tile_X14Y12_N1BEG;
	wire [7:0] Tile_X14Y12_N2BEG;
	wire [7:0] Tile_X14Y12_N2BEGb;
	wire [15:0] Tile_X14Y12_N4BEG;
	wire [15:0] Tile_X14Y12_NN4BEG;
	wire [0:0] Tile_X14Y12_Co;
	wire [3:0] Tile_X14Y12_E1BEG;
	wire [7:0] Tile_X14Y12_E2BEG;
	wire [7:0] Tile_X14Y12_E2BEGb;
	wire [15:0] Tile_X14Y12_EE4BEG;
	wire [11:0] Tile_X14Y12_E6BEG;
	wire [3:0] Tile_X14Y12_S1BEG;
	wire [7:0] Tile_X14Y12_S2BEG;
	wire [7:0] Tile_X14Y12_S2BEGb;
	wire [15:0] Tile_X14Y12_S4BEG;
	wire [15:0] Tile_X14Y12_SS4BEG;
	wire [3:0] Tile_X14Y12_W1BEG;
	wire [7:0] Tile_X14Y12_W2BEG;
	wire [7:0] Tile_X14Y12_W2BEGb;
	wire [15:0] Tile_X14Y12_WW4BEG;
	wire [11:0] Tile_X14Y12_W6BEG;
	wire [3:0] Tile_X15Y12_N1BEG;
	wire [7:0] Tile_X15Y12_N2BEG;
	wire [7:0] Tile_X15Y12_N2BEGb;
	wire [15:0] Tile_X15Y12_N4BEG;
	wire [3:0] Tile_X15Y12_S1BEG;
	wire [7:0] Tile_X15Y12_S2BEG;
	wire [7:0] Tile_X15Y12_S2BEGb;
	wire [15:0] Tile_X15Y12_S4BEG;
	wire [3:0] Tile_X15Y12_W1BEG;
	wire [7:0] Tile_X15Y12_W2BEG;
	wire [7:0] Tile_X15Y12_W2BEGb;
	wire [15:0] Tile_X15Y12_WW4BEG;
	wire [11:0] Tile_X15Y12_W6BEG;
	wire [3:0] Tile_X1Y13_N1BEG;
	wire [7:0] Tile_X1Y13_N2BEG;
	wire [7:0] Tile_X1Y13_N2BEGb;
	wire [15:0] Tile_X1Y13_N4BEG;
	wire [15:0] Tile_X1Y13_NN4BEG;
	wire [0:0] Tile_X1Y13_Co;
	wire [3:0] Tile_X2Y13_N1BEG;
	wire [7:0] Tile_X2Y13_N2BEG;
	wire [7:0] Tile_X2Y13_N2BEGb;
	wire [15:0] Tile_X2Y13_N4BEG;
	wire [15:0] Tile_X2Y13_NN4BEG;
	wire [3:0] Tile_X3Y13_N1BEG;
	wire [7:0] Tile_X3Y13_N2BEG;
	wire [7:0] Tile_X3Y13_N2BEGb;
	wire [15:0] Tile_X3Y13_N4BEG;
	wire [15:0] Tile_X3Y13_NN4BEG;
	wire [0:0] Tile_X3Y13_Co;
	wire [3:0] Tile_X4Y13_N1BEG;
	wire [7:0] Tile_X4Y13_N2BEG;
	wire [7:0] Tile_X4Y13_N2BEGb;
	wire [15:0] Tile_X4Y13_N4BEG;
	wire [15:0] Tile_X4Y13_NN4BEG;
	wire [0:0] Tile_X4Y13_Co;
	wire [3:0] Tile_X5Y13_N1BEG;
	wire [7:0] Tile_X5Y13_N2BEG;
	wire [7:0] Tile_X5Y13_N2BEGb;
	wire [15:0] Tile_X5Y13_N4BEG;
	wire [15:0] Tile_X5Y13_NN4BEG;
	wire [3:0] Tile_X6Y13_N1BEG;
	wire [7:0] Tile_X6Y13_N2BEG;
	wire [7:0] Tile_X6Y13_N2BEGb;
	wire [15:0] Tile_X6Y13_N4BEG;
	wire [15:0] Tile_X6Y13_NN4BEG;
	wire [0:0] Tile_X6Y13_Co;
	wire [3:0] Tile_X7Y13_N1BEG;
	wire [7:0] Tile_X7Y13_N2BEG;
	wire [7:0] Tile_X7Y13_N2BEGb;
	wire [15:0] Tile_X7Y13_N4BEG;
	wire [15:0] Tile_X7Y13_NN4BEG;
	wire [0:0] Tile_X7Y13_Co;
	wire [3:0] Tile_X8Y13_N1BEG;
	wire [7:0] Tile_X8Y13_N2BEG;
	wire [7:0] Tile_X8Y13_N2BEGb;
	wire [15:0] Tile_X8Y13_N4BEG;
	wire [15:0] Tile_X8Y13_NN4BEG;
	wire [0:0] Tile_X8Y13_Co;
	wire [3:0] Tile_X9Y13_N1BEG;
	wire [7:0] Tile_X9Y13_N2BEG;
	wire [7:0] Tile_X9Y13_N2BEGb;
	wire [15:0] Tile_X9Y13_N4BEG;
	wire [15:0] Tile_X9Y13_NN4BEG;
	wire [3:0] Tile_X10Y13_N1BEG;
	wire [7:0] Tile_X10Y13_N2BEG;
	wire [7:0] Tile_X10Y13_N2BEGb;
	wire [15:0] Tile_X10Y13_N4BEG;
	wire [15:0] Tile_X10Y13_NN4BEG;
	wire [0:0] Tile_X10Y13_Co;
	wire [3:0] Tile_X11Y13_N1BEG;
	wire [7:0] Tile_X11Y13_N2BEG;
	wire [7:0] Tile_X11Y13_N2BEGb;
	wire [15:0] Tile_X11Y13_N4BEG;
	wire [15:0] Tile_X11Y13_NN4BEG;
	wire [0:0] Tile_X11Y13_Co;
	wire [3:0] Tile_X12Y13_N1BEG;
	wire [7:0] Tile_X12Y13_N2BEG;
	wire [7:0] Tile_X12Y13_N2BEGb;
	wire [15:0] Tile_X12Y13_N4BEG;
	wire [15:0] Tile_X12Y13_NN4BEG;
	wire [0:0] Tile_X12Y13_Co;
	wire [3:0] Tile_X13Y13_N1BEG;
	wire [7:0] Tile_X13Y13_N2BEG;
	wire [7:0] Tile_X13Y13_N2BEGb;
	wire [15:0] Tile_X13Y13_N4BEG;
	wire [15:0] Tile_X13Y13_NN4BEG;
	wire [3:0] Tile_X14Y13_N1BEG;
	wire [7:0] Tile_X14Y13_N2BEG;
	wire [7:0] Tile_X14Y13_N2BEGb;
	wire [15:0] Tile_X14Y13_N4BEG;
	wire [15:0] Tile_X14Y13_NN4BEG;
	wire [0:0] Tile_X14Y13_Co;
	wire [3:0] Tile_X15Y13_N1BEG;
	wire [7:0] Tile_X15Y13_N2BEG;
	wire [7:0] Tile_X15Y13_N2BEGb;
	wire [15:0] Tile_X15Y13_N4BEG;

	assign Tile_Y1_FrameData = FrameData[(FrameBitsPerRow*(1+1))-1:FrameBitsPerRow*1];
	assign Tile_Y2_FrameData = FrameData[(FrameBitsPerRow*(2+1))-1:FrameBitsPerRow*2];
	assign Tile_Y3_FrameData = FrameData[(FrameBitsPerRow*(3+1))-1:FrameBitsPerRow*3];
	assign Tile_Y4_FrameData = FrameData[(FrameBitsPerRow*(4+1))-1:FrameBitsPerRow*4];
	assign Tile_Y5_FrameData = FrameData[(FrameBitsPerRow*(5+1))-1:FrameBitsPerRow*5];
	assign Tile_Y6_FrameData = FrameData[(FrameBitsPerRow*(6+1))-1:FrameBitsPerRow*6];
	assign Tile_Y7_FrameData = FrameData[(FrameBitsPerRow*(7+1))-1:FrameBitsPerRow*7];
	assign Tile_Y8_FrameData = FrameData[(FrameBitsPerRow*(8+1))-1:FrameBitsPerRow*8];
	assign Tile_Y9_FrameData = FrameData[(FrameBitsPerRow*(9+1))-1:FrameBitsPerRow*9];
	assign Tile_Y10_FrameData = FrameData[(FrameBitsPerRow*(10+1))-1:FrameBitsPerRow*10];
	assign Tile_Y11_FrameData = FrameData[(FrameBitsPerRow*(11+1))-1:FrameBitsPerRow*11];
	assign Tile_Y12_FrameData = FrameData[(FrameBitsPerRow*(12+1))-1:FrameBitsPerRow*12];
	assign Tile_X0_FrameStrobe = FrameStrobe[(MaxFramesPerCol*(0+1))-1:MaxFramesPerCol*0];
	assign Tile_X1_FrameStrobe = FrameStrobe[(MaxFramesPerCol*(1+1))-1:MaxFramesPerCol*1];
	assign Tile_X2_FrameStrobe = FrameStrobe[(MaxFramesPerCol*(2+1))-1:MaxFramesPerCol*2];
	assign Tile_X3_FrameStrobe = FrameStrobe[(MaxFramesPerCol*(3+1))-1:MaxFramesPerCol*3];
	assign Tile_X4_FrameStrobe = FrameStrobe[(MaxFramesPerCol*(4+1))-1:MaxFramesPerCol*4];
	assign Tile_X5_FrameStrobe = FrameStrobe[(MaxFramesPerCol*(5+1))-1:MaxFramesPerCol*5];
	assign Tile_X6_FrameStrobe = FrameStrobe[(MaxFramesPerCol*(6+1))-1:MaxFramesPerCol*6];
	assign Tile_X7_FrameStrobe = FrameStrobe[(MaxFramesPerCol*(7+1))-1:MaxFramesPerCol*7];
	assign Tile_X8_FrameStrobe = FrameStrobe[(MaxFramesPerCol*(8+1))-1:MaxFramesPerCol*8];
	assign Tile_X9_FrameStrobe = FrameStrobe[(MaxFramesPerCol*(9+1))-1:MaxFramesPerCol*9];
	assign Tile_X10_FrameStrobe = FrameStrobe[(MaxFramesPerCol*(10+1))-1:MaxFramesPerCol*10];
	assign Tile_X11_FrameStrobe = FrameStrobe[(MaxFramesPerCol*(11+1))-1:MaxFramesPerCol*11];
	assign Tile_X12_FrameStrobe = FrameStrobe[(MaxFramesPerCol*(12+1))-1:MaxFramesPerCol*12];
	assign Tile_X13_FrameStrobe = FrameStrobe[(MaxFramesPerCol*(13+1))-1:MaxFramesPerCol*13];
	assign Tile_X14_FrameStrobe = FrameStrobe[(MaxFramesPerCol*(14+1))-1:MaxFramesPerCol*14];
	assign Tile_X15_FrameStrobe = FrameStrobe[(MaxFramesPerCol*(15+1))-1:MaxFramesPerCol*15];

//tile instantiations

	N_term_DSP Tile_X5Y0_N_term_DSP (
	.N1END(Tile_X5Y1_N1BEG[3:0]),
	.N2MID(Tile_X5Y1_N2BEG[7:0]),
	.N2END(Tile_X5Y1_N2BEGb[7:0]),
	.N4END(Tile_X5Y1_N4BEG[15:0]),
	.NN4END(Tile_X5Y1_NN4BEG[15:0]),
	.S1BEG(Tile_X5Y0_S1BEG[3:0]),
	.S2BEG(Tile_X5Y0_S2BEG[7:0]),
	.S2BEGb(Tile_X5Y0_S2BEGb[7:0]),
	.S4BEG(Tile_X5Y0_S4BEG[15:0]),
	.SS4BEG(Tile_X5Y0_SS4BEG[15:0]),
	.UserCLK(Tile_X5Y1_UserCLKo),
	.UserCLKo(Tile_X5Y0_UserCLKo),
	.FrameStrobe(Tile_X5Y1_FrameStrobe_O),
	.FrameStrobe_O(Tile_X5Y0_FrameStrobe_O)
	);

	N_term_single Tile_X6Y0_N_term_single (
	.N1END(Tile_X6Y1_N1BEG[3:0]),
	.N2MID(Tile_X6Y1_N2BEG[7:0]),
	.N2END(Tile_X6Y1_N2BEGb[7:0]),
	.N4END(Tile_X6Y1_N4BEG[15:0]),
	.NN4END(Tile_X6Y1_NN4BEG[15:0]),
	.Ci(Tile_X6Y1_Co[0:0]),
	.S1BEG(Tile_X6Y0_S1BEG[3:0]),
	.S2BEG(Tile_X6Y0_S2BEG[7:0]),
	.S2BEGb(Tile_X6Y0_S2BEGb[7:0]),
	.S4BEG(Tile_X6Y0_S4BEG[15:0]),
	.SS4BEG(Tile_X6Y0_SS4BEG[15:0]),
	.UserCLK(Tile_X6Y1_UserCLKo),
	.UserCLKo(Tile_X6Y0_UserCLKo),
	.FrameStrobe(Tile_X6Y1_FrameStrobe_O),
	.FrameStrobe_O(Tile_X6Y0_FrameStrobe_O)
	);

	N_term_single Tile_X7Y0_N_term_single (
	.N1END(Tile_X7Y1_N1BEG[3:0]),
	.N2MID(Tile_X7Y1_N2BEG[7:0]),
	.N2END(Tile_X7Y1_N2BEGb[7:0]),
	.N4END(Tile_X7Y1_N4BEG[15:0]),
	.NN4END(Tile_X7Y1_NN4BEG[15:0]),
	.Ci(Tile_X7Y1_Co[0:0]),
	.S1BEG(Tile_X7Y0_S1BEG[3:0]),
	.S2BEG(Tile_X7Y0_S2BEG[7:0]),
	.S2BEGb(Tile_X7Y0_S2BEGb[7:0]),
	.S4BEG(Tile_X7Y0_S4BEG[15:0]),
	.SS4BEG(Tile_X7Y0_SS4BEG[15:0]),
	.UserCLK(Tile_X7Y1_UserCLKo),
	.UserCLKo(Tile_X7Y0_UserCLKo),
	.FrameStrobe(Tile_X7Y1_FrameStrobe_O),
	.FrameStrobe_O(Tile_X7Y0_FrameStrobe_O)
	);

	N_term_single Tile_X8Y0_N_term_single (
	.N1END(Tile_X8Y1_N1BEG[3:0]),
	.N2MID(Tile_X8Y1_N2BEG[7:0]),
	.N2END(Tile_X8Y1_N2BEGb[7:0]),
	.N4END(Tile_X8Y1_N4BEG[15:0]),
	.NN4END(Tile_X8Y1_NN4BEG[15:0]),
	.Ci(Tile_X8Y1_Co[0:0]),
	.S1BEG(Tile_X8Y0_S1BEG[3:0]),
	.S2BEG(Tile_X8Y0_S2BEG[7:0]),
	.S2BEGb(Tile_X8Y0_S2BEGb[7:0]),
	.S4BEG(Tile_X8Y0_S4BEG[15:0]),
	.SS4BEG(Tile_X8Y0_SS4BEG[15:0]),
	.UserCLK(Tile_X8Y1_UserCLKo),
	.UserCLKo(Tile_X8Y0_UserCLKo),
	.FrameStrobe(Tile_X8Y1_FrameStrobe_O),
	.FrameStrobe_O(Tile_X8Y0_FrameStrobe_O)
	);

	N_term_DSP Tile_X9Y0_N_term_DSP (
	.N1END(Tile_X9Y1_N1BEG[3:0]),
	.N2MID(Tile_X9Y1_N2BEG[7:0]),
	.N2END(Tile_X9Y1_N2BEGb[7:0]),
	.N4END(Tile_X9Y1_N4BEG[15:0]),
	.NN4END(Tile_X9Y1_NN4BEG[15:0]),
	.S1BEG(Tile_X9Y0_S1BEG[3:0]),
	.S2BEG(Tile_X9Y0_S2BEG[7:0]),
	.S2BEGb(Tile_X9Y0_S2BEGb[7:0]),
	.S4BEG(Tile_X9Y0_S4BEG[15:0]),
	.SS4BEG(Tile_X9Y0_SS4BEG[15:0]),
	.UserCLK(Tile_X9Y1_UserCLKo),
	.UserCLKo(Tile_X9Y0_UserCLKo),
	.FrameStrobe(Tile_X9Y1_FrameStrobe_O),
	.FrameStrobe_O(Tile_X9Y0_FrameStrobe_O)
	);

	N_term_single Tile_X10Y0_N_term_single (
	.N1END(Tile_X10Y1_N1BEG[3:0]),
	.N2MID(Tile_X10Y1_N2BEG[7:0]),
	.N2END(Tile_X10Y1_N2BEGb[7:0]),
	.N4END(Tile_X10Y1_N4BEG[15:0]),
	.NN4END(Tile_X10Y1_NN4BEG[15:0]),
	.Ci(Tile_X10Y1_Co[0:0]),
	.S1BEG(Tile_X10Y0_S1BEG[3:0]),
	.S2BEG(Tile_X10Y0_S2BEG[7:0]),
	.S2BEGb(Tile_X10Y0_S2BEGb[7:0]),
	.S4BEG(Tile_X10Y0_S4BEG[15:0]),
	.SS4BEG(Tile_X10Y0_SS4BEG[15:0]),
	.UserCLK(Tile_X10Y1_UserCLKo),
	.UserCLKo(Tile_X10Y0_UserCLKo),
	.FrameStrobe(Tile_X10Y1_FrameStrobe_O),
	.FrameStrobe_O(Tile_X10Y0_FrameStrobe_O)
	);

	W_CPU_IO Tile_X4Y1_W_CPU_IO (
	.W1END(Tile_X5Y1_W1BEG[3:0]),
	.W2MID(Tile_X5Y1_W2BEG[7:0]),
	.W2END(Tile_X5Y1_W2BEGb[7:0]),
	.WW4END(Tile_X5Y1_WW4BEG[15:0]),
	.W6END(Tile_X5Y1_W6BEG[11:0]),
	.E1BEG(Tile_X4Y1_E1BEG[3:0]),
	.E2BEG(Tile_X4Y1_E2BEG[7:0]),
	.E2BEGb(Tile_X4Y1_E2BEGb[7:0]),
	.EE4BEG(Tile_X4Y1_EE4BEG[15:0]),
	.E6BEG(Tile_X4Y1_E6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X4Y1_OPA_I0),
	.OPA_I1(Tile_X4Y1_OPA_I1),
	.OPA_I2(Tile_X4Y1_OPA_I2),
	.OPA_I3(Tile_X4Y1_OPA_I3),
	.UserCLK(Tile_X4Y2_UserCLKo),
	.OPB_I0(Tile_X4Y1_OPB_I0),
	.OPB_I1(Tile_X4Y1_OPB_I1),
	.OPB_I2(Tile_X4Y1_OPB_I2),
	.OPB_I3(Tile_X4Y1_OPB_I3),
	.RES0_O0(Tile_X4Y1_RES0_O0),
	.RES0_O1(Tile_X4Y1_RES0_O1),
	.RES0_O2(Tile_X4Y1_RES0_O2),
	.RES0_O3(Tile_X4Y1_RES0_O3),
	.RES1_O0(Tile_X4Y1_RES1_O0),
	.RES1_O1(Tile_X4Y1_RES1_O1),
	.RES1_O2(Tile_X4Y1_RES1_O2),
	.RES1_O3(Tile_X4Y1_RES1_O3),
	.RES2_O0(Tile_X4Y1_RES2_O0),
	.RES2_O1(Tile_X4Y1_RES2_O1),
	.RES2_O2(Tile_X4Y1_RES2_O2),
	.RES2_O3(Tile_X4Y1_RES2_O3),
	.UserCLKo(Tile_X4Y1_UserCLKo),
	.FrameData(Tile_Y1_FrameData), 
	.FrameData_O(Tile_X4Y1_FrameData_O), 
	.FrameStrobe(Tile_X4Y2_FrameStrobe_O),
	.FrameStrobe_O(Tile_X4Y1_FrameStrobe_O)
	);


	LUT4AB Tile_X6Y1_LUT4AB (
	.N1END(Tile_X6Y2_N1BEG[3:0]),
	.N2MID(Tile_X6Y2_N2BEG[7:0]),
	.N2END(Tile_X6Y2_N2BEGb[7:0]),
	.N4END(Tile_X6Y2_N4BEG[15:0]),
	.NN4END(Tile_X6Y2_NN4BEG[15:0]),
	.Ci(Tile_X6Y2_Co[0:0]),
	.E1END(Tile_X5Y1_E1BEG[3:0]),
	.E2MID(Tile_X5Y1_E2BEG[7:0]),
	.E2END(Tile_X5Y1_E2BEGb[7:0]),
	.EE4END(Tile_X5Y1_EE4BEG[15:0]),
	.E6END(Tile_X5Y1_E6BEG[11:0]),
	.S1END(Tile_X6Y0_S1BEG[3:0]),
	.S2MID(Tile_X6Y0_S2BEG[7:0]),
	.S2END(Tile_X6Y0_S2BEGb[7:0]),
	.S4END(Tile_X6Y0_S4BEG[15:0]),
	.SS4END(Tile_X6Y0_SS4BEG[15:0]),
	.W1END(Tile_X7Y1_W1BEG[3:0]),
	.W2MID(Tile_X7Y1_W2BEG[7:0]),
	.W2END(Tile_X7Y1_W2BEGb[7:0]),
	.WW4END(Tile_X7Y1_WW4BEG[15:0]),
	.W6END(Tile_X7Y1_W6BEG[11:0]),
	.N1BEG(Tile_X6Y1_N1BEG[3:0]),
	.N2BEG(Tile_X6Y1_N2BEG[7:0]),
	.N2BEGb(Tile_X6Y1_N2BEGb[7:0]),
	.N4BEG(Tile_X6Y1_N4BEG[15:0]),
	.NN4BEG(Tile_X6Y1_NN4BEG[15:0]),
	.Co(Tile_X6Y1_Co[0:0]),
	.E1BEG(Tile_X6Y1_E1BEG[3:0]),
	.E2BEG(Tile_X6Y1_E2BEG[7:0]),
	.E2BEGb(Tile_X6Y1_E2BEGb[7:0]),
	.EE4BEG(Tile_X6Y1_EE4BEG[15:0]),
	.E6BEG(Tile_X6Y1_E6BEG[11:0]),
	.S1BEG(Tile_X6Y1_S1BEG[3:0]),
	.S2BEG(Tile_X6Y1_S2BEG[7:0]),
	.S2BEGb(Tile_X6Y1_S2BEGb[7:0]),
	.S4BEG(Tile_X6Y1_S4BEG[15:0]),
	.SS4BEG(Tile_X6Y1_SS4BEG[15:0]),
	.W1BEG(Tile_X6Y1_W1BEG[3:0]),
	.W2BEG(Tile_X6Y1_W2BEG[7:0]),
	.W2BEGb(Tile_X6Y1_W2BEGb[7:0]),
	.WW4BEG(Tile_X6Y1_WW4BEG[15:0]),
	.W6BEG(Tile_X6Y1_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X6Y2_UserCLKo),
	.UserCLKo(Tile_X6Y1_UserCLKo),
	.FrameData(Tile_X5Y1_FrameData_O), 
	.FrameData_O(Tile_X6Y1_FrameData_O), 
	.FrameStrobe(Tile_X6Y2_FrameStrobe_O),
	.FrameStrobe_O(Tile_X6Y1_FrameStrobe_O)
	);

	LUT4AB Tile_X7Y1_LUT4AB (
	.N1END(Tile_X7Y2_N1BEG[3:0]),
	.N2MID(Tile_X7Y2_N2BEG[7:0]),
	.N2END(Tile_X7Y2_N2BEGb[7:0]),
	.N4END(Tile_X7Y2_N4BEG[15:0]),
	.NN4END(Tile_X7Y2_NN4BEG[15:0]),
	.Ci(Tile_X7Y2_Co[0:0]),
	.E1END(Tile_X6Y1_E1BEG[3:0]),
	.E2MID(Tile_X6Y1_E2BEG[7:0]),
	.E2END(Tile_X6Y1_E2BEGb[7:0]),
	.EE4END(Tile_X6Y1_EE4BEG[15:0]),
	.E6END(Tile_X6Y1_E6BEG[11:0]),
	.S1END(Tile_X7Y0_S1BEG[3:0]),
	.S2MID(Tile_X7Y0_S2BEG[7:0]),
	.S2END(Tile_X7Y0_S2BEGb[7:0]),
	.S4END(Tile_X7Y0_S4BEG[15:0]),
	.SS4END(Tile_X7Y0_SS4BEG[15:0]),
	.W1END(Tile_X8Y1_W1BEG[3:0]),
	.W2MID(Tile_X8Y1_W2BEG[7:0]),
	.W2END(Tile_X8Y1_W2BEGb[7:0]),
	.WW4END(Tile_X8Y1_WW4BEG[15:0]),
	.W6END(Tile_X8Y1_W6BEG[11:0]),
	.N1BEG(Tile_X7Y1_N1BEG[3:0]),
	.N2BEG(Tile_X7Y1_N2BEG[7:0]),
	.N2BEGb(Tile_X7Y1_N2BEGb[7:0]),
	.N4BEG(Tile_X7Y1_N4BEG[15:0]),
	.NN4BEG(Tile_X7Y1_NN4BEG[15:0]),
	.Co(Tile_X7Y1_Co[0:0]),
	.E1BEG(Tile_X7Y1_E1BEG[3:0]),
	.E2BEG(Tile_X7Y1_E2BEG[7:0]),
	.E2BEGb(Tile_X7Y1_E2BEGb[7:0]),
	.EE4BEG(Tile_X7Y1_EE4BEG[15:0]),
	.E6BEG(Tile_X7Y1_E6BEG[11:0]),
	.S1BEG(Tile_X7Y1_S1BEG[3:0]),
	.S2BEG(Tile_X7Y1_S2BEG[7:0]),
	.S2BEGb(Tile_X7Y1_S2BEGb[7:0]),
	.S4BEG(Tile_X7Y1_S4BEG[15:0]),
	.SS4BEG(Tile_X7Y1_SS4BEG[15:0]),
	.W1BEG(Tile_X7Y1_W1BEG[3:0]),
	.W2BEG(Tile_X7Y1_W2BEG[7:0]),
	.W2BEGb(Tile_X7Y1_W2BEGb[7:0]),
	.WW4BEG(Tile_X7Y1_WW4BEG[15:0]),
	.W6BEG(Tile_X7Y1_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X7Y2_UserCLKo),
	.UserCLKo(Tile_X7Y1_UserCLKo),
	.FrameData(Tile_X6Y1_FrameData_O), 
	.FrameData_O(Tile_X7Y1_FrameData_O), 
	.FrameStrobe(Tile_X7Y2_FrameStrobe_O),
	.FrameStrobe_O(Tile_X7Y1_FrameStrobe_O)
	);

	LUT4AB Tile_X8Y1_LUT4AB (
	.N1END(Tile_X8Y2_N1BEG[3:0]),
	.N2MID(Tile_X8Y2_N2BEG[7:0]),
	.N2END(Tile_X8Y2_N2BEGb[7:0]),
	.N4END(Tile_X8Y2_N4BEG[15:0]),
	.NN4END(Tile_X8Y2_NN4BEG[15:0]),
	.Ci(Tile_X8Y2_Co[0:0]),
	.E1END(Tile_X7Y1_E1BEG[3:0]),
	.E2MID(Tile_X7Y1_E2BEG[7:0]),
	.E2END(Tile_X7Y1_E2BEGb[7:0]),
	.EE4END(Tile_X7Y1_EE4BEG[15:0]),
	.E6END(Tile_X7Y1_E6BEG[11:0]),
	.S1END(Tile_X8Y0_S1BEG[3:0]),
	.S2MID(Tile_X8Y0_S2BEG[7:0]),
	.S2END(Tile_X8Y0_S2BEGb[7:0]),
	.S4END(Tile_X8Y0_S4BEG[15:0]),
	.SS4END(Tile_X8Y0_SS4BEG[15:0]),
	.W1END(Tile_X9Y1_W1BEG[3:0]),
	.W2MID(Tile_X9Y1_W2BEG[7:0]),
	.W2END(Tile_X9Y1_W2BEGb[7:0]),
	.WW4END(Tile_X9Y1_WW4BEG[15:0]),
	.W6END(Tile_X9Y1_W6BEG[11:0]),
	.N1BEG(Tile_X8Y1_N1BEG[3:0]),
	.N2BEG(Tile_X8Y1_N2BEG[7:0]),
	.N2BEGb(Tile_X8Y1_N2BEGb[7:0]),
	.N4BEG(Tile_X8Y1_N4BEG[15:0]),
	.NN4BEG(Tile_X8Y1_NN4BEG[15:0]),
	.Co(Tile_X8Y1_Co[0:0]),
	.E1BEG(Tile_X8Y1_E1BEG[3:0]),
	.E2BEG(Tile_X8Y1_E2BEG[7:0]),
	.E2BEGb(Tile_X8Y1_E2BEGb[7:0]),
	.EE4BEG(Tile_X8Y1_EE4BEG[15:0]),
	.E6BEG(Tile_X8Y1_E6BEG[11:0]),
	.S1BEG(Tile_X8Y1_S1BEG[3:0]),
	.S2BEG(Tile_X8Y1_S2BEG[7:0]),
	.S2BEGb(Tile_X8Y1_S2BEGb[7:0]),
	.S4BEG(Tile_X8Y1_S4BEG[15:0]),
	.SS4BEG(Tile_X8Y1_SS4BEG[15:0]),
	.W1BEG(Tile_X8Y1_W1BEG[3:0]),
	.W2BEG(Tile_X8Y1_W2BEG[7:0]),
	.W2BEGb(Tile_X8Y1_W2BEGb[7:0]),
	.WW4BEG(Tile_X8Y1_WW4BEG[15:0]),
	.W6BEG(Tile_X8Y1_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X8Y2_UserCLKo),
	.UserCLKo(Tile_X8Y1_UserCLKo),
	.FrameData(Tile_X7Y1_FrameData_O), 
	.FrameData_O(Tile_X8Y1_FrameData_O), 
	.FrameStrobe(Tile_X8Y2_FrameStrobe_O),
	.FrameStrobe_O(Tile_X8Y1_FrameStrobe_O)
	);


	LUT4AB Tile_X10Y1_LUT4AB (
	.N1END(Tile_X10Y2_N1BEG[3:0]),
	.N2MID(Tile_X10Y2_N2BEG[7:0]),
	.N2END(Tile_X10Y2_N2BEGb[7:0]),
	.N4END(Tile_X10Y2_N4BEG[15:0]),
	.NN4END(Tile_X10Y2_NN4BEG[15:0]),
	.Ci(Tile_X10Y2_Co[0:0]),
	.E1END(Tile_X9Y1_E1BEG[3:0]),
	.E2MID(Tile_X9Y1_E2BEG[7:0]),
	.E2END(Tile_X9Y1_E2BEGb[7:0]),
	.EE4END(Tile_X9Y1_EE4BEG[15:0]),
	.E6END(Tile_X9Y1_E6BEG[11:0]),
	.S1END(Tile_X10Y0_S1BEG[3:0]),
	.S2MID(Tile_X10Y0_S2BEG[7:0]),
	.S2END(Tile_X10Y0_S2BEGb[7:0]),
	.S4END(Tile_X10Y0_S4BEG[15:0]),
	.SS4END(Tile_X10Y0_SS4BEG[15:0]),
	.W1END(Tile_X11Y1_W1BEG[3:0]),
	.W2MID(Tile_X11Y1_W2BEG[7:0]),
	.W2END(Tile_X11Y1_W2BEGb[7:0]),
	.WW4END(Tile_X11Y1_WW4BEG[15:0]),
	.W6END(Tile_X11Y1_W6BEG[11:0]),
	.N1BEG(Tile_X10Y1_N1BEG[3:0]),
	.N2BEG(Tile_X10Y1_N2BEG[7:0]),
	.N2BEGb(Tile_X10Y1_N2BEGb[7:0]),
	.N4BEG(Tile_X10Y1_N4BEG[15:0]),
	.NN4BEG(Tile_X10Y1_NN4BEG[15:0]),
	.Co(Tile_X10Y1_Co[0:0]),
	.E1BEG(Tile_X10Y1_E1BEG[3:0]),
	.E2BEG(Tile_X10Y1_E2BEG[7:0]),
	.E2BEGb(Tile_X10Y1_E2BEGb[7:0]),
	.EE4BEG(Tile_X10Y1_EE4BEG[15:0]),
	.E6BEG(Tile_X10Y1_E6BEG[11:0]),
	.S1BEG(Tile_X10Y1_S1BEG[3:0]),
	.S2BEG(Tile_X10Y1_S2BEG[7:0]),
	.S2BEGb(Tile_X10Y1_S2BEGb[7:0]),
	.S4BEG(Tile_X10Y1_S4BEG[15:0]),
	.SS4BEG(Tile_X10Y1_SS4BEG[15:0]),
	.W1BEG(Tile_X10Y1_W1BEG[3:0]),
	.W2BEG(Tile_X10Y1_W2BEG[7:0]),
	.W2BEGb(Tile_X10Y1_W2BEGb[7:0]),
	.WW4BEG(Tile_X10Y1_WW4BEG[15:0]),
	.W6BEG(Tile_X10Y1_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X10Y2_UserCLKo),
	.UserCLKo(Tile_X10Y1_UserCLKo),
	.FrameData(Tile_X9Y1_FrameData_O), 
	.FrameData_O(Tile_X10Y1_FrameData_O), 
	.FrameStrobe(Tile_X10Y2_FrameStrobe_O),
	.FrameStrobe_O(Tile_X10Y1_FrameStrobe_O)
	);

	E_CPU_IO Tile_X11Y1_E_CPU_IO (
	.E1END(Tile_X10Y1_E1BEG[3:0]),
	.E2MID(Tile_X10Y1_E2BEG[7:0]),
	.E2END(Tile_X10Y1_E2BEGb[7:0]),
	.EE4END(Tile_X10Y1_EE4BEG[15:0]),
	.E6END(Tile_X10Y1_E6BEG[11:0]),
	.W1BEG(Tile_X11Y1_W1BEG[3:0]),
	.W2BEG(Tile_X11Y1_W2BEG[7:0]),
	.W2BEGb(Tile_X11Y1_W2BEGb[7:0]),
	.WW4BEG(Tile_X11Y1_WW4BEG[15:0]),
	.W6BEG(Tile_X11Y1_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X11Y1_OPA_I0),
	.OPA_I1(Tile_X11Y1_OPA_I1),
	.OPA_I2(Tile_X11Y1_OPA_I2),
	.OPA_I3(Tile_X11Y1_OPA_I3),
	.UserCLK(Tile_X11Y2_UserCLKo),
	.OPB_I0(Tile_X11Y1_OPB_I0),
	.OPB_I1(Tile_X11Y1_OPB_I1),
	.OPB_I2(Tile_X11Y1_OPB_I2),
	.OPB_I3(Tile_X11Y1_OPB_I3),
	.RES0_O0(Tile_X11Y1_RES0_O0),
	.RES0_O1(Tile_X11Y1_RES0_O1),
	.RES0_O2(Tile_X11Y1_RES0_O2),
	.RES0_O3(Tile_X11Y1_RES0_O3),
	.RES1_O0(Tile_X11Y1_RES1_O0),
	.RES1_O1(Tile_X11Y1_RES1_O1),
	.RES1_O2(Tile_X11Y1_RES1_O2),
	.RES1_O3(Tile_X11Y1_RES1_O3),
	.RES2_O0(Tile_X11Y1_RES2_O0),
	.RES2_O1(Tile_X11Y1_RES2_O1),
	.RES2_O2(Tile_X11Y1_RES2_O2),
	.RES2_O3(Tile_X11Y1_RES2_O3),
	.UserCLKo(Tile_X11Y1_UserCLKo),
	.FrameData(Tile_X10Y1_FrameData_O), 
	.FrameData_O(Tile_X11Y1_FrameData_O), 
	.FrameStrobe(Tile_X11Y2_FrameStrobe_O),
	.FrameStrobe_O(Tile_X11Y1_FrameStrobe_O)
	);

	W_CPU_IO Tile_X4Y2_W_CPU_IO (
	.W1END(Tile_X5Y2_W1BEG[3:0]),
	.W2MID(Tile_X5Y2_W2BEG[7:0]),
	.W2END(Tile_X5Y2_W2BEGb[7:0]),
	.WW4END(Tile_X5Y2_WW4BEG[15:0]),
	.W6END(Tile_X5Y2_W6BEG[11:0]),
	.E1BEG(Tile_X4Y2_E1BEG[3:0]),
	.E2BEG(Tile_X4Y2_E2BEG[7:0]),
	.E2BEGb(Tile_X4Y2_E2BEGb[7:0]),
	.EE4BEG(Tile_X4Y2_EE4BEG[15:0]),
	.E6BEG(Tile_X4Y2_E6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X4Y2_OPA_I0),
	.OPA_I1(Tile_X4Y2_OPA_I1),
	.OPA_I2(Tile_X4Y2_OPA_I2),
	.OPA_I3(Tile_X4Y2_OPA_I3),
	.UserCLK(Tile_X4Y3_UserCLKo),
	.OPB_I0(Tile_X4Y2_OPB_I0),
	.OPB_I1(Tile_X4Y2_OPB_I1),
	.OPB_I2(Tile_X4Y2_OPB_I2),
	.OPB_I3(Tile_X4Y2_OPB_I3),
	.RES0_O0(Tile_X4Y2_RES0_O0),
	.RES0_O1(Tile_X4Y2_RES0_O1),
	.RES0_O2(Tile_X4Y2_RES0_O2),
	.RES0_O3(Tile_X4Y2_RES0_O3),
	.RES1_O0(Tile_X4Y2_RES1_O0),
	.RES1_O1(Tile_X4Y2_RES1_O1),
	.RES1_O2(Tile_X4Y2_RES1_O2),
	.RES1_O3(Tile_X4Y2_RES1_O3),
	.RES2_O0(Tile_X4Y2_RES2_O0),
	.RES2_O1(Tile_X4Y2_RES2_O1),
	.RES2_O2(Tile_X4Y2_RES2_O2),
	.RES2_O3(Tile_X4Y2_RES2_O3),
	.UserCLKo(Tile_X4Y2_UserCLKo),
	.FrameData(Tile_Y2_FrameData), 
	.FrameData_O(Tile_X4Y2_FrameData_O), 
	.FrameStrobe(Tile_X4Y3_FrameStrobe_O),
	.FrameStrobe_O(Tile_X4Y2_FrameStrobe_O)
	);


	LUT4AB Tile_X6Y2_LUT4AB (
	.N1END(Tile_X6Y3_N1BEG[3:0]),
	.N2MID(Tile_X6Y3_N2BEG[7:0]),
	.N2END(Tile_X6Y3_N2BEGb[7:0]),
	.N4END(Tile_X6Y3_N4BEG[15:0]),
	.NN4END(Tile_X6Y3_NN4BEG[15:0]),
	.Ci(Tile_X6Y3_Co[0:0]),
	.E1END(Tile_X5Y2_E1BEG[3:0]),
	.E2MID(Tile_X5Y2_E2BEG[7:0]),
	.E2END(Tile_X5Y2_E2BEGb[7:0]),
	.EE4END(Tile_X5Y2_EE4BEG[15:0]),
	.E6END(Tile_X5Y2_E6BEG[11:0]),
	.S1END(Tile_X6Y1_S1BEG[3:0]),
	.S2MID(Tile_X6Y1_S2BEG[7:0]),
	.S2END(Tile_X6Y1_S2BEGb[7:0]),
	.S4END(Tile_X6Y1_S4BEG[15:0]),
	.SS4END(Tile_X6Y1_SS4BEG[15:0]),
	.W1END(Tile_X7Y2_W1BEG[3:0]),
	.W2MID(Tile_X7Y2_W2BEG[7:0]),
	.W2END(Tile_X7Y2_W2BEGb[7:0]),
	.WW4END(Tile_X7Y2_WW4BEG[15:0]),
	.W6END(Tile_X7Y2_W6BEG[11:0]),
	.N1BEG(Tile_X6Y2_N1BEG[3:0]),
	.N2BEG(Tile_X6Y2_N2BEG[7:0]),
	.N2BEGb(Tile_X6Y2_N2BEGb[7:0]),
	.N4BEG(Tile_X6Y2_N4BEG[15:0]),
	.NN4BEG(Tile_X6Y2_NN4BEG[15:0]),
	.Co(Tile_X6Y2_Co[0:0]),
	.E1BEG(Tile_X6Y2_E1BEG[3:0]),
	.E2BEG(Tile_X6Y2_E2BEG[7:0]),
	.E2BEGb(Tile_X6Y2_E2BEGb[7:0]),
	.EE4BEG(Tile_X6Y2_EE4BEG[15:0]),
	.E6BEG(Tile_X6Y2_E6BEG[11:0]),
	.S1BEG(Tile_X6Y2_S1BEG[3:0]),
	.S2BEG(Tile_X6Y2_S2BEG[7:0]),
	.S2BEGb(Tile_X6Y2_S2BEGb[7:0]),
	.S4BEG(Tile_X6Y2_S4BEG[15:0]),
	.SS4BEG(Tile_X6Y2_SS4BEG[15:0]),
	.W1BEG(Tile_X6Y2_W1BEG[3:0]),
	.W2BEG(Tile_X6Y2_W2BEG[7:0]),
	.W2BEGb(Tile_X6Y2_W2BEGb[7:0]),
	.WW4BEG(Tile_X6Y2_WW4BEG[15:0]),
	.W6BEG(Tile_X6Y2_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X6Y3_UserCLKo),
	.UserCLKo(Tile_X6Y2_UserCLKo),
	.FrameData(Tile_X5Y2_FrameData_O), 
	.FrameData_O(Tile_X6Y2_FrameData_O), 
	.FrameStrobe(Tile_X6Y3_FrameStrobe_O),
	.FrameStrobe_O(Tile_X6Y2_FrameStrobe_O)
	);

	LUT4AB Tile_X7Y2_LUT4AB (
	.N1END(Tile_X7Y3_N1BEG[3:0]),
	.N2MID(Tile_X7Y3_N2BEG[7:0]),
	.N2END(Tile_X7Y3_N2BEGb[7:0]),
	.N4END(Tile_X7Y3_N4BEG[15:0]),
	.NN4END(Tile_X7Y3_NN4BEG[15:0]),
	.Ci(Tile_X7Y3_Co[0:0]),
	.E1END(Tile_X6Y2_E1BEG[3:0]),
	.E2MID(Tile_X6Y2_E2BEG[7:0]),
	.E2END(Tile_X6Y2_E2BEGb[7:0]),
	.EE4END(Tile_X6Y2_EE4BEG[15:0]),
	.E6END(Tile_X6Y2_E6BEG[11:0]),
	.S1END(Tile_X7Y1_S1BEG[3:0]),
	.S2MID(Tile_X7Y1_S2BEG[7:0]),
	.S2END(Tile_X7Y1_S2BEGb[7:0]),
	.S4END(Tile_X7Y1_S4BEG[15:0]),
	.SS4END(Tile_X7Y1_SS4BEG[15:0]),
	.W1END(Tile_X8Y2_W1BEG[3:0]),
	.W2MID(Tile_X8Y2_W2BEG[7:0]),
	.W2END(Tile_X8Y2_W2BEGb[7:0]),
	.WW4END(Tile_X8Y2_WW4BEG[15:0]),
	.W6END(Tile_X8Y2_W6BEG[11:0]),
	.N1BEG(Tile_X7Y2_N1BEG[3:0]),
	.N2BEG(Tile_X7Y2_N2BEG[7:0]),
	.N2BEGb(Tile_X7Y2_N2BEGb[7:0]),
	.N4BEG(Tile_X7Y2_N4BEG[15:0]),
	.NN4BEG(Tile_X7Y2_NN4BEG[15:0]),
	.Co(Tile_X7Y2_Co[0:0]),
	.E1BEG(Tile_X7Y2_E1BEG[3:0]),
	.E2BEG(Tile_X7Y2_E2BEG[7:0]),
	.E2BEGb(Tile_X7Y2_E2BEGb[7:0]),
	.EE4BEG(Tile_X7Y2_EE4BEG[15:0]),
	.E6BEG(Tile_X7Y2_E6BEG[11:0]),
	.S1BEG(Tile_X7Y2_S1BEG[3:0]),
	.S2BEG(Tile_X7Y2_S2BEG[7:0]),
	.S2BEGb(Tile_X7Y2_S2BEGb[7:0]),
	.S4BEG(Tile_X7Y2_S4BEG[15:0]),
	.SS4BEG(Tile_X7Y2_SS4BEG[15:0]),
	.W1BEG(Tile_X7Y2_W1BEG[3:0]),
	.W2BEG(Tile_X7Y2_W2BEG[7:0]),
	.W2BEGb(Tile_X7Y2_W2BEGb[7:0]),
	.WW4BEG(Tile_X7Y2_WW4BEG[15:0]),
	.W6BEG(Tile_X7Y2_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X7Y3_UserCLKo),
	.UserCLKo(Tile_X7Y2_UserCLKo),
	.FrameData(Tile_X6Y2_FrameData_O), 
	.FrameData_O(Tile_X7Y2_FrameData_O), 
	.FrameStrobe(Tile_X7Y3_FrameStrobe_O),
	.FrameStrobe_O(Tile_X7Y2_FrameStrobe_O)
	);

	LUT4AB Tile_X8Y2_LUT4AB (
	.N1END(Tile_X8Y3_N1BEG[3:0]),
	.N2MID(Tile_X8Y3_N2BEG[7:0]),
	.N2END(Tile_X8Y3_N2BEGb[7:0]),
	.N4END(Tile_X8Y3_N4BEG[15:0]),
	.NN4END(Tile_X8Y3_NN4BEG[15:0]),
	.Ci(Tile_X8Y3_Co[0:0]),
	.E1END(Tile_X7Y2_E1BEG[3:0]),
	.E2MID(Tile_X7Y2_E2BEG[7:0]),
	.E2END(Tile_X7Y2_E2BEGb[7:0]),
	.EE4END(Tile_X7Y2_EE4BEG[15:0]),
	.E6END(Tile_X7Y2_E6BEG[11:0]),
	.S1END(Tile_X8Y1_S1BEG[3:0]),
	.S2MID(Tile_X8Y1_S2BEG[7:0]),
	.S2END(Tile_X8Y1_S2BEGb[7:0]),
	.S4END(Tile_X8Y1_S4BEG[15:0]),
	.SS4END(Tile_X8Y1_SS4BEG[15:0]),
	.W1END(Tile_X9Y2_W1BEG[3:0]),
	.W2MID(Tile_X9Y2_W2BEG[7:0]),
	.W2END(Tile_X9Y2_W2BEGb[7:0]),
	.WW4END(Tile_X9Y2_WW4BEG[15:0]),
	.W6END(Tile_X9Y2_W6BEG[11:0]),
	.N1BEG(Tile_X8Y2_N1BEG[3:0]),
	.N2BEG(Tile_X8Y2_N2BEG[7:0]),
	.N2BEGb(Tile_X8Y2_N2BEGb[7:0]),
	.N4BEG(Tile_X8Y2_N4BEG[15:0]),
	.NN4BEG(Tile_X8Y2_NN4BEG[15:0]),
	.Co(Tile_X8Y2_Co[0:0]),
	.E1BEG(Tile_X8Y2_E1BEG[3:0]),
	.E2BEG(Tile_X8Y2_E2BEG[7:0]),
	.E2BEGb(Tile_X8Y2_E2BEGb[7:0]),
	.EE4BEG(Tile_X8Y2_EE4BEG[15:0]),
	.E6BEG(Tile_X8Y2_E6BEG[11:0]),
	.S1BEG(Tile_X8Y2_S1BEG[3:0]),
	.S2BEG(Tile_X8Y2_S2BEG[7:0]),
	.S2BEGb(Tile_X8Y2_S2BEGb[7:0]),
	.S4BEG(Tile_X8Y2_S4BEG[15:0]),
	.SS4BEG(Tile_X8Y2_SS4BEG[15:0]),
	.W1BEG(Tile_X8Y2_W1BEG[3:0]),
	.W2BEG(Tile_X8Y2_W2BEG[7:0]),
	.W2BEGb(Tile_X8Y2_W2BEGb[7:0]),
	.WW4BEG(Tile_X8Y2_WW4BEG[15:0]),
	.W6BEG(Tile_X8Y2_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X8Y3_UserCLKo),
	.UserCLKo(Tile_X8Y2_UserCLKo),
	.FrameData(Tile_X7Y2_FrameData_O), 
	.FrameData_O(Tile_X8Y2_FrameData_O), 
	.FrameStrobe(Tile_X8Y3_FrameStrobe_O),
	.FrameStrobe_O(Tile_X8Y2_FrameStrobe_O)
	);


	LUT4AB Tile_X10Y2_LUT4AB (
	.N1END(Tile_X10Y3_N1BEG[3:0]),
	.N2MID(Tile_X10Y3_N2BEG[7:0]),
	.N2END(Tile_X10Y3_N2BEGb[7:0]),
	.N4END(Tile_X10Y3_N4BEG[15:0]),
	.NN4END(Tile_X10Y3_NN4BEG[15:0]),
	.Ci(Tile_X10Y3_Co[0:0]),
	.E1END(Tile_X9Y2_E1BEG[3:0]),
	.E2MID(Tile_X9Y2_E2BEG[7:0]),
	.E2END(Tile_X9Y2_E2BEGb[7:0]),
	.EE4END(Tile_X9Y2_EE4BEG[15:0]),
	.E6END(Tile_X9Y2_E6BEG[11:0]),
	.S1END(Tile_X10Y1_S1BEG[3:0]),
	.S2MID(Tile_X10Y1_S2BEG[7:0]),
	.S2END(Tile_X10Y1_S2BEGb[7:0]),
	.S4END(Tile_X10Y1_S4BEG[15:0]),
	.SS4END(Tile_X10Y1_SS4BEG[15:0]),
	.W1END(Tile_X11Y2_W1BEG[3:0]),
	.W2MID(Tile_X11Y2_W2BEG[7:0]),
	.W2END(Tile_X11Y2_W2BEGb[7:0]),
	.WW4END(Tile_X11Y2_WW4BEG[15:0]),
	.W6END(Tile_X11Y2_W6BEG[11:0]),
	.N1BEG(Tile_X10Y2_N1BEG[3:0]),
	.N2BEG(Tile_X10Y2_N2BEG[7:0]),
	.N2BEGb(Tile_X10Y2_N2BEGb[7:0]),
	.N4BEG(Tile_X10Y2_N4BEG[15:0]),
	.NN4BEG(Tile_X10Y2_NN4BEG[15:0]),
	.Co(Tile_X10Y2_Co[0:0]),
	.E1BEG(Tile_X10Y2_E1BEG[3:0]),
	.E2BEG(Tile_X10Y2_E2BEG[7:0]),
	.E2BEGb(Tile_X10Y2_E2BEGb[7:0]),
	.EE4BEG(Tile_X10Y2_EE4BEG[15:0]),
	.E6BEG(Tile_X10Y2_E6BEG[11:0]),
	.S1BEG(Tile_X10Y2_S1BEG[3:0]),
	.S2BEG(Tile_X10Y2_S2BEG[7:0]),
	.S2BEGb(Tile_X10Y2_S2BEGb[7:0]),
	.S4BEG(Tile_X10Y2_S4BEG[15:0]),
	.SS4BEG(Tile_X10Y2_SS4BEG[15:0]),
	.W1BEG(Tile_X10Y2_W1BEG[3:0]),
	.W2BEG(Tile_X10Y2_W2BEG[7:0]),
	.W2BEGb(Tile_X10Y2_W2BEGb[7:0]),
	.WW4BEG(Tile_X10Y2_WW4BEG[15:0]),
	.W6BEG(Tile_X10Y2_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X10Y3_UserCLKo),
	.UserCLKo(Tile_X10Y2_UserCLKo),
	.FrameData(Tile_X9Y2_FrameData_O), 
	.FrameData_O(Tile_X10Y2_FrameData_O), 
	.FrameStrobe(Tile_X10Y3_FrameStrobe_O),
	.FrameStrobe_O(Tile_X10Y2_FrameStrobe_O)
	);

	E_CPU_IO Tile_X11Y2_E_CPU_IO (
	.E1END(Tile_X10Y2_E1BEG[3:0]),
	.E2MID(Tile_X10Y2_E2BEG[7:0]),
	.E2END(Tile_X10Y2_E2BEGb[7:0]),
	.EE4END(Tile_X10Y2_EE4BEG[15:0]),
	.E6END(Tile_X10Y2_E6BEG[11:0]),
	.W1BEG(Tile_X11Y2_W1BEG[3:0]),
	.W2BEG(Tile_X11Y2_W2BEG[7:0]),
	.W2BEGb(Tile_X11Y2_W2BEGb[7:0]),
	.WW4BEG(Tile_X11Y2_WW4BEG[15:0]),
	.W6BEG(Tile_X11Y2_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X11Y2_OPA_I0),
	.OPA_I1(Tile_X11Y2_OPA_I1),
	.OPA_I2(Tile_X11Y2_OPA_I2),
	.OPA_I3(Tile_X11Y2_OPA_I3),
	.UserCLK(Tile_X11Y3_UserCLKo),
	.OPB_I0(Tile_X11Y2_OPB_I0),
	.OPB_I1(Tile_X11Y2_OPB_I1),
	.OPB_I2(Tile_X11Y2_OPB_I2),
	.OPB_I3(Tile_X11Y2_OPB_I3),
	.RES0_O0(Tile_X11Y2_RES0_O0),
	.RES0_O1(Tile_X11Y2_RES0_O1),
	.RES0_O2(Tile_X11Y2_RES0_O2),
	.RES0_O3(Tile_X11Y2_RES0_O3),
	.RES1_O0(Tile_X11Y2_RES1_O0),
	.RES1_O1(Tile_X11Y2_RES1_O1),
	.RES1_O2(Tile_X11Y2_RES1_O2),
	.RES1_O3(Tile_X11Y2_RES1_O3),
	.RES2_O0(Tile_X11Y2_RES2_O0),
	.RES2_O1(Tile_X11Y2_RES2_O1),
	.RES2_O2(Tile_X11Y2_RES2_O2),
	.RES2_O3(Tile_X11Y2_RES2_O3),
	.UserCLKo(Tile_X11Y2_UserCLKo),
	.FrameData(Tile_X10Y2_FrameData_O), 
	.FrameData_O(Tile_X11Y2_FrameData_O), 
	.FrameStrobe(Tile_X11Y3_FrameStrobe_O),
	.FrameStrobe_O(Tile_X11Y2_FrameStrobe_O)
	);

	W_CPU_IO Tile_X4Y3_W_CPU_IO (
	.W1END(Tile_X5Y3_W1BEG[3:0]),
	.W2MID(Tile_X5Y3_W2BEG[7:0]),
	.W2END(Tile_X5Y3_W2BEGb[7:0]),
	.WW4END(Tile_X5Y3_WW4BEG[15:0]),
	.W6END(Tile_X5Y3_W6BEG[11:0]),
	.E1BEG(Tile_X4Y3_E1BEG[3:0]),
	.E2BEG(Tile_X4Y3_E2BEG[7:0]),
	.E2BEGb(Tile_X4Y3_E2BEGb[7:0]),
	.EE4BEG(Tile_X4Y3_EE4BEG[15:0]),
	.E6BEG(Tile_X4Y3_E6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X4Y3_OPA_I0),
	.OPA_I1(Tile_X4Y3_OPA_I1),
	.OPA_I2(Tile_X4Y3_OPA_I2),
	.OPA_I3(Tile_X4Y3_OPA_I3),
	.UserCLK(Tile_X4Y4_UserCLKo),
	.OPB_I0(Tile_X4Y3_OPB_I0),
	.OPB_I1(Tile_X4Y3_OPB_I1),
	.OPB_I2(Tile_X4Y3_OPB_I2),
	.OPB_I3(Tile_X4Y3_OPB_I3),
	.RES0_O0(Tile_X4Y3_RES0_O0),
	.RES0_O1(Tile_X4Y3_RES0_O1),
	.RES0_O2(Tile_X4Y3_RES0_O2),
	.RES0_O3(Tile_X4Y3_RES0_O3),
	.RES1_O0(Tile_X4Y3_RES1_O0),
	.RES1_O1(Tile_X4Y3_RES1_O1),
	.RES1_O2(Tile_X4Y3_RES1_O2),
	.RES1_O3(Tile_X4Y3_RES1_O3),
	.RES2_O0(Tile_X4Y3_RES2_O0),
	.RES2_O1(Tile_X4Y3_RES2_O1),
	.RES2_O2(Tile_X4Y3_RES2_O2),
	.RES2_O3(Tile_X4Y3_RES2_O3),
	.UserCLKo(Tile_X4Y3_UserCLKo),
	.FrameData(Tile_Y3_FrameData), 
	.FrameData_O(Tile_X4Y3_FrameData_O), 
	.FrameStrobe(Tile_X4Y4_FrameStrobe_O),
	.FrameStrobe_O(Tile_X4Y3_FrameStrobe_O)
	);


	LUT4AB Tile_X6Y3_LUT4AB (
	.N1END(Tile_X6Y4_N1BEG[3:0]),
	.N2MID(Tile_X6Y4_N2BEG[7:0]),
	.N2END(Tile_X6Y4_N2BEGb[7:0]),
	.N4END(Tile_X6Y4_N4BEG[15:0]),
	.NN4END(Tile_X6Y4_NN4BEG[15:0]),
	.Ci(Tile_X6Y4_Co[0:0]),
	.E1END(Tile_X5Y3_E1BEG[3:0]),
	.E2MID(Tile_X5Y3_E2BEG[7:0]),
	.E2END(Tile_X5Y3_E2BEGb[7:0]),
	.EE4END(Tile_X5Y3_EE4BEG[15:0]),
	.E6END(Tile_X5Y3_E6BEG[11:0]),
	.S1END(Tile_X6Y2_S1BEG[3:0]),
	.S2MID(Tile_X6Y2_S2BEG[7:0]),
	.S2END(Tile_X6Y2_S2BEGb[7:0]),
	.S4END(Tile_X6Y2_S4BEG[15:0]),
	.SS4END(Tile_X6Y2_SS4BEG[15:0]),
	.W1END(Tile_X7Y3_W1BEG[3:0]),
	.W2MID(Tile_X7Y3_W2BEG[7:0]),
	.W2END(Tile_X7Y3_W2BEGb[7:0]),
	.WW4END(Tile_X7Y3_WW4BEG[15:0]),
	.W6END(Tile_X7Y3_W6BEG[11:0]),
	.N1BEG(Tile_X6Y3_N1BEG[3:0]),
	.N2BEG(Tile_X6Y3_N2BEG[7:0]),
	.N2BEGb(Tile_X6Y3_N2BEGb[7:0]),
	.N4BEG(Tile_X6Y3_N4BEG[15:0]),
	.NN4BEG(Tile_X6Y3_NN4BEG[15:0]),
	.Co(Tile_X6Y3_Co[0:0]),
	.E1BEG(Tile_X6Y3_E1BEG[3:0]),
	.E2BEG(Tile_X6Y3_E2BEG[7:0]),
	.E2BEGb(Tile_X6Y3_E2BEGb[7:0]),
	.EE4BEG(Tile_X6Y3_EE4BEG[15:0]),
	.E6BEG(Tile_X6Y3_E6BEG[11:0]),
	.S1BEG(Tile_X6Y3_S1BEG[3:0]),
	.S2BEG(Tile_X6Y3_S2BEG[7:0]),
	.S2BEGb(Tile_X6Y3_S2BEGb[7:0]),
	.S4BEG(Tile_X6Y3_S4BEG[15:0]),
	.SS4BEG(Tile_X6Y3_SS4BEG[15:0]),
	.W1BEG(Tile_X6Y3_W1BEG[3:0]),
	.W2BEG(Tile_X6Y3_W2BEG[7:0]),
	.W2BEGb(Tile_X6Y3_W2BEGb[7:0]),
	.WW4BEG(Tile_X6Y3_WW4BEG[15:0]),
	.W6BEG(Tile_X6Y3_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X6Y4_UserCLKo),
	.UserCLKo(Tile_X6Y3_UserCLKo),
	.FrameData(Tile_X5Y3_FrameData_O), 
	.FrameData_O(Tile_X6Y3_FrameData_O), 
	.FrameStrobe(Tile_X6Y4_FrameStrobe_O),
	.FrameStrobe_O(Tile_X6Y3_FrameStrobe_O)
	);

	LUT4AB Tile_X7Y3_LUT4AB (
	.N1END(Tile_X7Y4_N1BEG[3:0]),
	.N2MID(Tile_X7Y4_N2BEG[7:0]),
	.N2END(Tile_X7Y4_N2BEGb[7:0]),
	.N4END(Tile_X7Y4_N4BEG[15:0]),
	.NN4END(Tile_X7Y4_NN4BEG[15:0]),
	.Ci(Tile_X7Y4_Co[0:0]),
	.E1END(Tile_X6Y3_E1BEG[3:0]),
	.E2MID(Tile_X6Y3_E2BEG[7:0]),
	.E2END(Tile_X6Y3_E2BEGb[7:0]),
	.EE4END(Tile_X6Y3_EE4BEG[15:0]),
	.E6END(Tile_X6Y3_E6BEG[11:0]),
	.S1END(Tile_X7Y2_S1BEG[3:0]),
	.S2MID(Tile_X7Y2_S2BEG[7:0]),
	.S2END(Tile_X7Y2_S2BEGb[7:0]),
	.S4END(Tile_X7Y2_S4BEG[15:0]),
	.SS4END(Tile_X7Y2_SS4BEG[15:0]),
	.W1END(Tile_X8Y3_W1BEG[3:0]),
	.W2MID(Tile_X8Y3_W2BEG[7:0]),
	.W2END(Tile_X8Y3_W2BEGb[7:0]),
	.WW4END(Tile_X8Y3_WW4BEG[15:0]),
	.W6END(Tile_X8Y3_W6BEG[11:0]),
	.N1BEG(Tile_X7Y3_N1BEG[3:0]),
	.N2BEG(Tile_X7Y3_N2BEG[7:0]),
	.N2BEGb(Tile_X7Y3_N2BEGb[7:0]),
	.N4BEG(Tile_X7Y3_N4BEG[15:0]),
	.NN4BEG(Tile_X7Y3_NN4BEG[15:0]),
	.Co(Tile_X7Y3_Co[0:0]),
	.E1BEG(Tile_X7Y3_E1BEG[3:0]),
	.E2BEG(Tile_X7Y3_E2BEG[7:0]),
	.E2BEGb(Tile_X7Y3_E2BEGb[7:0]),
	.EE4BEG(Tile_X7Y3_EE4BEG[15:0]),
	.E6BEG(Tile_X7Y3_E6BEG[11:0]),
	.S1BEG(Tile_X7Y3_S1BEG[3:0]),
	.S2BEG(Tile_X7Y3_S2BEG[7:0]),
	.S2BEGb(Tile_X7Y3_S2BEGb[7:0]),
	.S4BEG(Tile_X7Y3_S4BEG[15:0]),
	.SS4BEG(Tile_X7Y3_SS4BEG[15:0]),
	.W1BEG(Tile_X7Y3_W1BEG[3:0]),
	.W2BEG(Tile_X7Y3_W2BEG[7:0]),
	.W2BEGb(Tile_X7Y3_W2BEGb[7:0]),
	.WW4BEG(Tile_X7Y3_WW4BEG[15:0]),
	.W6BEG(Tile_X7Y3_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X7Y4_UserCLKo),
	.UserCLKo(Tile_X7Y3_UserCLKo),
	.FrameData(Tile_X6Y3_FrameData_O), 
	.FrameData_O(Tile_X7Y3_FrameData_O), 
	.FrameStrobe(Tile_X7Y4_FrameStrobe_O),
	.FrameStrobe_O(Tile_X7Y3_FrameStrobe_O)
	);

	LUT4AB Tile_X8Y3_LUT4AB (
	.N1END(Tile_X8Y4_N1BEG[3:0]),
	.N2MID(Tile_X8Y4_N2BEG[7:0]),
	.N2END(Tile_X8Y4_N2BEGb[7:0]),
	.N4END(Tile_X8Y4_N4BEG[15:0]),
	.NN4END(Tile_X8Y4_NN4BEG[15:0]),
	.Ci(Tile_X8Y4_Co[0:0]),
	.E1END(Tile_X7Y3_E1BEG[3:0]),
	.E2MID(Tile_X7Y3_E2BEG[7:0]),
	.E2END(Tile_X7Y3_E2BEGb[7:0]),
	.EE4END(Tile_X7Y3_EE4BEG[15:0]),
	.E6END(Tile_X7Y3_E6BEG[11:0]),
	.S1END(Tile_X8Y2_S1BEG[3:0]),
	.S2MID(Tile_X8Y2_S2BEG[7:0]),
	.S2END(Tile_X8Y2_S2BEGb[7:0]),
	.S4END(Tile_X8Y2_S4BEG[15:0]),
	.SS4END(Tile_X8Y2_SS4BEG[15:0]),
	.W1END(Tile_X9Y3_W1BEG[3:0]),
	.W2MID(Tile_X9Y3_W2BEG[7:0]),
	.W2END(Tile_X9Y3_W2BEGb[7:0]),
	.WW4END(Tile_X9Y3_WW4BEG[15:0]),
	.W6END(Tile_X9Y3_W6BEG[11:0]),
	.N1BEG(Tile_X8Y3_N1BEG[3:0]),
	.N2BEG(Tile_X8Y3_N2BEG[7:0]),
	.N2BEGb(Tile_X8Y3_N2BEGb[7:0]),
	.N4BEG(Tile_X8Y3_N4BEG[15:0]),
	.NN4BEG(Tile_X8Y3_NN4BEG[15:0]),
	.Co(Tile_X8Y3_Co[0:0]),
	.E1BEG(Tile_X8Y3_E1BEG[3:0]),
	.E2BEG(Tile_X8Y3_E2BEG[7:0]),
	.E2BEGb(Tile_X8Y3_E2BEGb[7:0]),
	.EE4BEG(Tile_X8Y3_EE4BEG[15:0]),
	.E6BEG(Tile_X8Y3_E6BEG[11:0]),
	.S1BEG(Tile_X8Y3_S1BEG[3:0]),
	.S2BEG(Tile_X8Y3_S2BEG[7:0]),
	.S2BEGb(Tile_X8Y3_S2BEGb[7:0]),
	.S4BEG(Tile_X8Y3_S4BEG[15:0]),
	.SS4BEG(Tile_X8Y3_SS4BEG[15:0]),
	.W1BEG(Tile_X8Y3_W1BEG[3:0]),
	.W2BEG(Tile_X8Y3_W2BEG[7:0]),
	.W2BEGb(Tile_X8Y3_W2BEGb[7:0]),
	.WW4BEG(Tile_X8Y3_WW4BEG[15:0]),
	.W6BEG(Tile_X8Y3_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X8Y4_UserCLKo),
	.UserCLKo(Tile_X8Y3_UserCLKo),
	.FrameData(Tile_X7Y3_FrameData_O), 
	.FrameData_O(Tile_X8Y3_FrameData_O), 
	.FrameStrobe(Tile_X8Y4_FrameStrobe_O),
	.FrameStrobe_O(Tile_X8Y3_FrameStrobe_O)
	);


	LUT4AB Tile_X10Y3_LUT4AB (
	.N1END(Tile_X10Y4_N1BEG[3:0]),
	.N2MID(Tile_X10Y4_N2BEG[7:0]),
	.N2END(Tile_X10Y4_N2BEGb[7:0]),
	.N4END(Tile_X10Y4_N4BEG[15:0]),
	.NN4END(Tile_X10Y4_NN4BEG[15:0]),
	.Ci(Tile_X10Y4_Co[0:0]),
	.E1END(Tile_X9Y3_E1BEG[3:0]),
	.E2MID(Tile_X9Y3_E2BEG[7:0]),
	.E2END(Tile_X9Y3_E2BEGb[7:0]),
	.EE4END(Tile_X9Y3_EE4BEG[15:0]),
	.E6END(Tile_X9Y3_E6BEG[11:0]),
	.S1END(Tile_X10Y2_S1BEG[3:0]),
	.S2MID(Tile_X10Y2_S2BEG[7:0]),
	.S2END(Tile_X10Y2_S2BEGb[7:0]),
	.S4END(Tile_X10Y2_S4BEG[15:0]),
	.SS4END(Tile_X10Y2_SS4BEG[15:0]),
	.W1END(Tile_X11Y3_W1BEG[3:0]),
	.W2MID(Tile_X11Y3_W2BEG[7:0]),
	.W2END(Tile_X11Y3_W2BEGb[7:0]),
	.WW4END(Tile_X11Y3_WW4BEG[15:0]),
	.W6END(Tile_X11Y3_W6BEG[11:0]),
	.N1BEG(Tile_X10Y3_N1BEG[3:0]),
	.N2BEG(Tile_X10Y3_N2BEG[7:0]),
	.N2BEGb(Tile_X10Y3_N2BEGb[7:0]),
	.N4BEG(Tile_X10Y3_N4BEG[15:0]),
	.NN4BEG(Tile_X10Y3_NN4BEG[15:0]),
	.Co(Tile_X10Y3_Co[0:0]),
	.E1BEG(Tile_X10Y3_E1BEG[3:0]),
	.E2BEG(Tile_X10Y3_E2BEG[7:0]),
	.E2BEGb(Tile_X10Y3_E2BEGb[7:0]),
	.EE4BEG(Tile_X10Y3_EE4BEG[15:0]),
	.E6BEG(Tile_X10Y3_E6BEG[11:0]),
	.S1BEG(Tile_X10Y3_S1BEG[3:0]),
	.S2BEG(Tile_X10Y3_S2BEG[7:0]),
	.S2BEGb(Tile_X10Y3_S2BEGb[7:0]),
	.S4BEG(Tile_X10Y3_S4BEG[15:0]),
	.SS4BEG(Tile_X10Y3_SS4BEG[15:0]),
	.W1BEG(Tile_X10Y3_W1BEG[3:0]),
	.W2BEG(Tile_X10Y3_W2BEG[7:0]),
	.W2BEGb(Tile_X10Y3_W2BEGb[7:0]),
	.WW4BEG(Tile_X10Y3_WW4BEG[15:0]),
	.W6BEG(Tile_X10Y3_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X10Y4_UserCLKo),
	.UserCLKo(Tile_X10Y3_UserCLKo),
	.FrameData(Tile_X9Y3_FrameData_O), 
	.FrameData_O(Tile_X10Y3_FrameData_O), 
	.FrameStrobe(Tile_X10Y4_FrameStrobe_O),
	.FrameStrobe_O(Tile_X10Y3_FrameStrobe_O)
	);

	E_CPU_IO Tile_X11Y3_E_CPU_IO (
	.E1END(Tile_X10Y3_E1BEG[3:0]),
	.E2MID(Tile_X10Y3_E2BEG[7:0]),
	.E2END(Tile_X10Y3_E2BEGb[7:0]),
	.EE4END(Tile_X10Y3_EE4BEG[15:0]),
	.E6END(Tile_X10Y3_E6BEG[11:0]),
	.W1BEG(Tile_X11Y3_W1BEG[3:0]),
	.W2BEG(Tile_X11Y3_W2BEG[7:0]),
	.W2BEGb(Tile_X11Y3_W2BEGb[7:0]),
	.WW4BEG(Tile_X11Y3_WW4BEG[15:0]),
	.W6BEG(Tile_X11Y3_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X11Y3_OPA_I0),
	.OPA_I1(Tile_X11Y3_OPA_I1),
	.OPA_I2(Tile_X11Y3_OPA_I2),
	.OPA_I3(Tile_X11Y3_OPA_I3),
	.UserCLK(Tile_X11Y4_UserCLKo),
	.OPB_I0(Tile_X11Y3_OPB_I0),
	.OPB_I1(Tile_X11Y3_OPB_I1),
	.OPB_I2(Tile_X11Y3_OPB_I2),
	.OPB_I3(Tile_X11Y3_OPB_I3),
	.RES0_O0(Tile_X11Y3_RES0_O0),
	.RES0_O1(Tile_X11Y3_RES0_O1),
	.RES0_O2(Tile_X11Y3_RES0_O2),
	.RES0_O3(Tile_X11Y3_RES0_O3),
	.RES1_O0(Tile_X11Y3_RES1_O0),
	.RES1_O1(Tile_X11Y3_RES1_O1),
	.RES1_O2(Tile_X11Y3_RES1_O2),
	.RES1_O3(Tile_X11Y3_RES1_O3),
	.RES2_O0(Tile_X11Y3_RES2_O0),
	.RES2_O1(Tile_X11Y3_RES2_O1),
	.RES2_O2(Tile_X11Y3_RES2_O2),
	.RES2_O3(Tile_X11Y3_RES2_O3),
	.UserCLKo(Tile_X11Y3_UserCLKo),
	.FrameData(Tile_X10Y3_FrameData_O), 
	.FrameData_O(Tile_X11Y3_FrameData_O), 
	.FrameStrobe(Tile_X11Y4_FrameStrobe_O),
	.FrameStrobe_O(Tile_X11Y3_FrameStrobe_O)
	);

	W_CPU_IO Tile_X4Y4_W_CPU_IO (
	.W1END(Tile_X5Y4_W1BEG[3:0]),
	.W2MID(Tile_X5Y4_W2BEG[7:0]),
	.W2END(Tile_X5Y4_W2BEGb[7:0]),
	.WW4END(Tile_X5Y4_WW4BEG[15:0]),
	.W6END(Tile_X5Y4_W6BEG[11:0]),
	.E1BEG(Tile_X4Y4_E1BEG[3:0]),
	.E2BEG(Tile_X4Y4_E2BEG[7:0]),
	.E2BEGb(Tile_X4Y4_E2BEGb[7:0]),
	.EE4BEG(Tile_X4Y4_EE4BEG[15:0]),
	.E6BEG(Tile_X4Y4_E6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X4Y4_OPA_I0),
	.OPA_I1(Tile_X4Y4_OPA_I1),
	.OPA_I2(Tile_X4Y4_OPA_I2),
	.OPA_I3(Tile_X4Y4_OPA_I3),
	.UserCLK(Tile_X4Y5_UserCLKo),
	.OPB_I0(Tile_X4Y4_OPB_I0),
	.OPB_I1(Tile_X4Y4_OPB_I1),
	.OPB_I2(Tile_X4Y4_OPB_I2),
	.OPB_I3(Tile_X4Y4_OPB_I3),
	.RES0_O0(Tile_X4Y4_RES0_O0),
	.RES0_O1(Tile_X4Y4_RES0_O1),
	.RES0_O2(Tile_X4Y4_RES0_O2),
	.RES0_O3(Tile_X4Y4_RES0_O3),
	.RES1_O0(Tile_X4Y4_RES1_O0),
	.RES1_O1(Tile_X4Y4_RES1_O1),
	.RES1_O2(Tile_X4Y4_RES1_O2),
	.RES1_O3(Tile_X4Y4_RES1_O3),
	.RES2_O0(Tile_X4Y4_RES2_O0),
	.RES2_O1(Tile_X4Y4_RES2_O1),
	.RES2_O2(Tile_X4Y4_RES2_O2),
	.RES2_O3(Tile_X4Y4_RES2_O3),
	.UserCLKo(Tile_X4Y4_UserCLKo),
	.FrameData(Tile_Y4_FrameData), 
	.FrameData_O(Tile_X4Y4_FrameData_O), 
	.FrameStrobe(Tile_X4Y5_FrameStrobe_O),
	.FrameStrobe_O(Tile_X4Y4_FrameStrobe_O)
	);


	LUT4AB Tile_X6Y4_LUT4AB (
	.N1END(Tile_X6Y5_N1BEG[3:0]),
	.N2MID(Tile_X6Y5_N2BEG[7:0]),
	.N2END(Tile_X6Y5_N2BEGb[7:0]),
	.N4END(Tile_X6Y5_N4BEG[15:0]),
	.NN4END(Tile_X6Y5_NN4BEG[15:0]),
	.Ci(Tile_X6Y5_Co[0:0]),
	.E1END(Tile_X5Y4_E1BEG[3:0]),
	.E2MID(Tile_X5Y4_E2BEG[7:0]),
	.E2END(Tile_X5Y4_E2BEGb[7:0]),
	.EE4END(Tile_X5Y4_EE4BEG[15:0]),
	.E6END(Tile_X5Y4_E6BEG[11:0]),
	.S1END(Tile_X6Y3_S1BEG[3:0]),
	.S2MID(Tile_X6Y3_S2BEG[7:0]),
	.S2END(Tile_X6Y3_S2BEGb[7:0]),
	.S4END(Tile_X6Y3_S4BEG[15:0]),
	.SS4END(Tile_X6Y3_SS4BEG[15:0]),
	.W1END(Tile_X7Y4_W1BEG[3:0]),
	.W2MID(Tile_X7Y4_W2BEG[7:0]),
	.W2END(Tile_X7Y4_W2BEGb[7:0]),
	.WW4END(Tile_X7Y4_WW4BEG[15:0]),
	.W6END(Tile_X7Y4_W6BEG[11:0]),
	.N1BEG(Tile_X6Y4_N1BEG[3:0]),
	.N2BEG(Tile_X6Y4_N2BEG[7:0]),
	.N2BEGb(Tile_X6Y4_N2BEGb[7:0]),
	.N4BEG(Tile_X6Y4_N4BEG[15:0]),
	.NN4BEG(Tile_X6Y4_NN4BEG[15:0]),
	.Co(Tile_X6Y4_Co[0:0]),
	.E1BEG(Tile_X6Y4_E1BEG[3:0]),
	.E2BEG(Tile_X6Y4_E2BEG[7:0]),
	.E2BEGb(Tile_X6Y4_E2BEGb[7:0]),
	.EE4BEG(Tile_X6Y4_EE4BEG[15:0]),
	.E6BEG(Tile_X6Y4_E6BEG[11:0]),
	.S1BEG(Tile_X6Y4_S1BEG[3:0]),
	.S2BEG(Tile_X6Y4_S2BEG[7:0]),
	.S2BEGb(Tile_X6Y4_S2BEGb[7:0]),
	.S4BEG(Tile_X6Y4_S4BEG[15:0]),
	.SS4BEG(Tile_X6Y4_SS4BEG[15:0]),
	.W1BEG(Tile_X6Y4_W1BEG[3:0]),
	.W2BEG(Tile_X6Y4_W2BEG[7:0]),
	.W2BEGb(Tile_X6Y4_W2BEGb[7:0]),
	.WW4BEG(Tile_X6Y4_WW4BEG[15:0]),
	.W6BEG(Tile_X6Y4_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X6Y5_UserCLKo),
	.UserCLKo(Tile_X6Y4_UserCLKo),
	.FrameData(Tile_X5Y4_FrameData_O), 
	.FrameData_O(Tile_X6Y4_FrameData_O), 
	.FrameStrobe(Tile_X6Y5_FrameStrobe_O),
	.FrameStrobe_O(Tile_X6Y4_FrameStrobe_O)
	);

	LUT4AB Tile_X7Y4_LUT4AB (
	.N1END(Tile_X7Y5_N1BEG[3:0]),
	.N2MID(Tile_X7Y5_N2BEG[7:0]),
	.N2END(Tile_X7Y5_N2BEGb[7:0]),
	.N4END(Tile_X7Y5_N4BEG[15:0]),
	.NN4END(Tile_X7Y5_NN4BEG[15:0]),
	.Ci(Tile_X7Y5_Co[0:0]),
	.E1END(Tile_X6Y4_E1BEG[3:0]),
	.E2MID(Tile_X6Y4_E2BEG[7:0]),
	.E2END(Tile_X6Y4_E2BEGb[7:0]),
	.EE4END(Tile_X6Y4_EE4BEG[15:0]),
	.E6END(Tile_X6Y4_E6BEG[11:0]),
	.S1END(Tile_X7Y3_S1BEG[3:0]),
	.S2MID(Tile_X7Y3_S2BEG[7:0]),
	.S2END(Tile_X7Y3_S2BEGb[7:0]),
	.S4END(Tile_X7Y3_S4BEG[15:0]),
	.SS4END(Tile_X7Y3_SS4BEG[15:0]),
	.W1END(Tile_X8Y4_W1BEG[3:0]),
	.W2MID(Tile_X8Y4_W2BEG[7:0]),
	.W2END(Tile_X8Y4_W2BEGb[7:0]),
	.WW4END(Tile_X8Y4_WW4BEG[15:0]),
	.W6END(Tile_X8Y4_W6BEG[11:0]),
	.N1BEG(Tile_X7Y4_N1BEG[3:0]),
	.N2BEG(Tile_X7Y4_N2BEG[7:0]),
	.N2BEGb(Tile_X7Y4_N2BEGb[7:0]),
	.N4BEG(Tile_X7Y4_N4BEG[15:0]),
	.NN4BEG(Tile_X7Y4_NN4BEG[15:0]),
	.Co(Tile_X7Y4_Co[0:0]),
	.E1BEG(Tile_X7Y4_E1BEG[3:0]),
	.E2BEG(Tile_X7Y4_E2BEG[7:0]),
	.E2BEGb(Tile_X7Y4_E2BEGb[7:0]),
	.EE4BEG(Tile_X7Y4_EE4BEG[15:0]),
	.E6BEG(Tile_X7Y4_E6BEG[11:0]),
	.S1BEG(Tile_X7Y4_S1BEG[3:0]),
	.S2BEG(Tile_X7Y4_S2BEG[7:0]),
	.S2BEGb(Tile_X7Y4_S2BEGb[7:0]),
	.S4BEG(Tile_X7Y4_S4BEG[15:0]),
	.SS4BEG(Tile_X7Y4_SS4BEG[15:0]),
	.W1BEG(Tile_X7Y4_W1BEG[3:0]),
	.W2BEG(Tile_X7Y4_W2BEG[7:0]),
	.W2BEGb(Tile_X7Y4_W2BEGb[7:0]),
	.WW4BEG(Tile_X7Y4_WW4BEG[15:0]),
	.W6BEG(Tile_X7Y4_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X7Y5_UserCLKo),
	.UserCLKo(Tile_X7Y4_UserCLKo),
	.FrameData(Tile_X6Y4_FrameData_O), 
	.FrameData_O(Tile_X7Y4_FrameData_O), 
	.FrameStrobe(Tile_X7Y5_FrameStrobe_O),
	.FrameStrobe_O(Tile_X7Y4_FrameStrobe_O)
	);

	LUT4AB Tile_X8Y4_LUT4AB (
	.N1END(Tile_X8Y5_N1BEG[3:0]),
	.N2MID(Tile_X8Y5_N2BEG[7:0]),
	.N2END(Tile_X8Y5_N2BEGb[7:0]),
	.N4END(Tile_X8Y5_N4BEG[15:0]),
	.NN4END(Tile_X8Y5_NN4BEG[15:0]),
	.Ci(Tile_X8Y5_Co[0:0]),
	.E1END(Tile_X7Y4_E1BEG[3:0]),
	.E2MID(Tile_X7Y4_E2BEG[7:0]),
	.E2END(Tile_X7Y4_E2BEGb[7:0]),
	.EE4END(Tile_X7Y4_EE4BEG[15:0]),
	.E6END(Tile_X7Y4_E6BEG[11:0]),
	.S1END(Tile_X8Y3_S1BEG[3:0]),
	.S2MID(Tile_X8Y3_S2BEG[7:0]),
	.S2END(Tile_X8Y3_S2BEGb[7:0]),
	.S4END(Tile_X8Y3_S4BEG[15:0]),
	.SS4END(Tile_X8Y3_SS4BEG[15:0]),
	.W1END(Tile_X9Y4_W1BEG[3:0]),
	.W2MID(Tile_X9Y4_W2BEG[7:0]),
	.W2END(Tile_X9Y4_W2BEGb[7:0]),
	.WW4END(Tile_X9Y4_WW4BEG[15:0]),
	.W6END(Tile_X9Y4_W6BEG[11:0]),
	.N1BEG(Tile_X8Y4_N1BEG[3:0]),
	.N2BEG(Tile_X8Y4_N2BEG[7:0]),
	.N2BEGb(Tile_X8Y4_N2BEGb[7:0]),
	.N4BEG(Tile_X8Y4_N4BEG[15:0]),
	.NN4BEG(Tile_X8Y4_NN4BEG[15:0]),
	.Co(Tile_X8Y4_Co[0:0]),
	.E1BEG(Tile_X8Y4_E1BEG[3:0]),
	.E2BEG(Tile_X8Y4_E2BEG[7:0]),
	.E2BEGb(Tile_X8Y4_E2BEGb[7:0]),
	.EE4BEG(Tile_X8Y4_EE4BEG[15:0]),
	.E6BEG(Tile_X8Y4_E6BEG[11:0]),
	.S1BEG(Tile_X8Y4_S1BEG[3:0]),
	.S2BEG(Tile_X8Y4_S2BEG[7:0]),
	.S2BEGb(Tile_X8Y4_S2BEGb[7:0]),
	.S4BEG(Tile_X8Y4_S4BEG[15:0]),
	.SS4BEG(Tile_X8Y4_SS4BEG[15:0]),
	.W1BEG(Tile_X8Y4_W1BEG[3:0]),
	.W2BEG(Tile_X8Y4_W2BEG[7:0]),
	.W2BEGb(Tile_X8Y4_W2BEGb[7:0]),
	.WW4BEG(Tile_X8Y4_WW4BEG[15:0]),
	.W6BEG(Tile_X8Y4_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X8Y5_UserCLKo),
	.UserCLKo(Tile_X8Y4_UserCLKo),
	.FrameData(Tile_X7Y4_FrameData_O), 
	.FrameData_O(Tile_X8Y4_FrameData_O), 
	.FrameStrobe(Tile_X8Y5_FrameStrobe_O),
	.FrameStrobe_O(Tile_X8Y4_FrameStrobe_O)
	);


	LUT4AB Tile_X10Y4_LUT4AB (
	.N1END(Tile_X10Y5_N1BEG[3:0]),
	.N2MID(Tile_X10Y5_N2BEG[7:0]),
	.N2END(Tile_X10Y5_N2BEGb[7:0]),
	.N4END(Tile_X10Y5_N4BEG[15:0]),
	.NN4END(Tile_X10Y5_NN4BEG[15:0]),
	.Ci(Tile_X10Y5_Co[0:0]),
	.E1END(Tile_X9Y4_E1BEG[3:0]),
	.E2MID(Tile_X9Y4_E2BEG[7:0]),
	.E2END(Tile_X9Y4_E2BEGb[7:0]),
	.EE4END(Tile_X9Y4_EE4BEG[15:0]),
	.E6END(Tile_X9Y4_E6BEG[11:0]),
	.S1END(Tile_X10Y3_S1BEG[3:0]),
	.S2MID(Tile_X10Y3_S2BEG[7:0]),
	.S2END(Tile_X10Y3_S2BEGb[7:0]),
	.S4END(Tile_X10Y3_S4BEG[15:0]),
	.SS4END(Tile_X10Y3_SS4BEG[15:0]),
	.W1END(Tile_X11Y4_W1BEG[3:0]),
	.W2MID(Tile_X11Y4_W2BEG[7:0]),
	.W2END(Tile_X11Y4_W2BEGb[7:0]),
	.WW4END(Tile_X11Y4_WW4BEG[15:0]),
	.W6END(Tile_X11Y4_W6BEG[11:0]),
	.N1BEG(Tile_X10Y4_N1BEG[3:0]),
	.N2BEG(Tile_X10Y4_N2BEG[7:0]),
	.N2BEGb(Tile_X10Y4_N2BEGb[7:0]),
	.N4BEG(Tile_X10Y4_N4BEG[15:0]),
	.NN4BEG(Tile_X10Y4_NN4BEG[15:0]),
	.Co(Tile_X10Y4_Co[0:0]),
	.E1BEG(Tile_X10Y4_E1BEG[3:0]),
	.E2BEG(Tile_X10Y4_E2BEG[7:0]),
	.E2BEGb(Tile_X10Y4_E2BEGb[7:0]),
	.EE4BEG(Tile_X10Y4_EE4BEG[15:0]),
	.E6BEG(Tile_X10Y4_E6BEG[11:0]),
	.S1BEG(Tile_X10Y4_S1BEG[3:0]),
	.S2BEG(Tile_X10Y4_S2BEG[7:0]),
	.S2BEGb(Tile_X10Y4_S2BEGb[7:0]),
	.S4BEG(Tile_X10Y4_S4BEG[15:0]),
	.SS4BEG(Tile_X10Y4_SS4BEG[15:0]),
	.W1BEG(Tile_X10Y4_W1BEG[3:0]),
	.W2BEG(Tile_X10Y4_W2BEG[7:0]),
	.W2BEGb(Tile_X10Y4_W2BEGb[7:0]),
	.WW4BEG(Tile_X10Y4_WW4BEG[15:0]),
	.W6BEG(Tile_X10Y4_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X10Y5_UserCLKo),
	.UserCLKo(Tile_X10Y4_UserCLKo),
	.FrameData(Tile_X9Y4_FrameData_O), 
	.FrameData_O(Tile_X10Y4_FrameData_O), 
	.FrameStrobe(Tile_X10Y5_FrameStrobe_O),
	.FrameStrobe_O(Tile_X10Y4_FrameStrobe_O)
	);

	E_CPU_IO Tile_X11Y4_E_CPU_IO (
	.E1END(Tile_X10Y4_E1BEG[3:0]),
	.E2MID(Tile_X10Y4_E2BEG[7:0]),
	.E2END(Tile_X10Y4_E2BEGb[7:0]),
	.EE4END(Tile_X10Y4_EE4BEG[15:0]),
	.E6END(Tile_X10Y4_E6BEG[11:0]),
	.W1BEG(Tile_X11Y4_W1BEG[3:0]),
	.W2BEG(Tile_X11Y4_W2BEG[7:0]),
	.W2BEGb(Tile_X11Y4_W2BEGb[7:0]),
	.WW4BEG(Tile_X11Y4_WW4BEG[15:0]),
	.W6BEG(Tile_X11Y4_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X11Y4_OPA_I0),
	.OPA_I1(Tile_X11Y4_OPA_I1),
	.OPA_I2(Tile_X11Y4_OPA_I2),
	.OPA_I3(Tile_X11Y4_OPA_I3),
	.UserCLK(Tile_X11Y5_UserCLKo),
	.OPB_I0(Tile_X11Y4_OPB_I0),
	.OPB_I1(Tile_X11Y4_OPB_I1),
	.OPB_I2(Tile_X11Y4_OPB_I2),
	.OPB_I3(Tile_X11Y4_OPB_I3),
	.RES0_O0(Tile_X11Y4_RES0_O0),
	.RES0_O1(Tile_X11Y4_RES0_O1),
	.RES0_O2(Tile_X11Y4_RES0_O2),
	.RES0_O3(Tile_X11Y4_RES0_O3),
	.RES1_O0(Tile_X11Y4_RES1_O0),
	.RES1_O1(Tile_X11Y4_RES1_O1),
	.RES1_O2(Tile_X11Y4_RES1_O2),
	.RES1_O3(Tile_X11Y4_RES1_O3),
	.RES2_O0(Tile_X11Y4_RES2_O0),
	.RES2_O1(Tile_X11Y4_RES2_O1),
	.RES2_O2(Tile_X11Y4_RES2_O2),
	.RES2_O3(Tile_X11Y4_RES2_O3),
	.UserCLKo(Tile_X11Y4_UserCLKo),
	.FrameData(Tile_X10Y4_FrameData_O), 
	.FrameData_O(Tile_X11Y4_FrameData_O), 
	.FrameStrobe(Tile_X11Y5_FrameStrobe_O),
	.FrameStrobe_O(Tile_X11Y4_FrameStrobe_O)
	);

	W_CPU_IO Tile_X4Y5_W_CPU_IO (
	.W1END(Tile_X5Y5_W1BEG[3:0]),
	.W2MID(Tile_X5Y5_W2BEG[7:0]),
	.W2END(Tile_X5Y5_W2BEGb[7:0]),
	.WW4END(Tile_X5Y5_WW4BEG[15:0]),
	.W6END(Tile_X5Y5_W6BEG[11:0]),
	.E1BEG(Tile_X4Y5_E1BEG[3:0]),
	.E2BEG(Tile_X4Y5_E2BEG[7:0]),
	.E2BEGb(Tile_X4Y5_E2BEGb[7:0]),
	.EE4BEG(Tile_X4Y5_EE4BEG[15:0]),
	.E6BEG(Tile_X4Y5_E6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X4Y5_OPA_I0),
	.OPA_I1(Tile_X4Y5_OPA_I1),
	.OPA_I2(Tile_X4Y5_OPA_I2),
	.OPA_I3(Tile_X4Y5_OPA_I3),
	.UserCLK(Tile_X4Y6_UserCLKo),
	.OPB_I0(Tile_X4Y5_OPB_I0),
	.OPB_I1(Tile_X4Y5_OPB_I1),
	.OPB_I2(Tile_X4Y5_OPB_I2),
	.OPB_I3(Tile_X4Y5_OPB_I3),
	.RES0_O0(Tile_X4Y5_RES0_O0),
	.RES0_O1(Tile_X4Y5_RES0_O1),
	.RES0_O2(Tile_X4Y5_RES0_O2),
	.RES0_O3(Tile_X4Y5_RES0_O3),
	.RES1_O0(Tile_X4Y5_RES1_O0),
	.RES1_O1(Tile_X4Y5_RES1_O1),
	.RES1_O2(Tile_X4Y5_RES1_O2),
	.RES1_O3(Tile_X4Y5_RES1_O3),
	.RES2_O0(Tile_X4Y5_RES2_O0),
	.RES2_O1(Tile_X4Y5_RES2_O1),
	.RES2_O2(Tile_X4Y5_RES2_O2),
	.RES2_O3(Tile_X4Y5_RES2_O3),
	.UserCLKo(Tile_X4Y5_UserCLKo),
	.FrameData(Tile_Y5_FrameData), 
	.FrameData_O(Tile_X4Y5_FrameData_O), 
	.FrameStrobe(Tile_X4Y6_FrameStrobe_O),
	.FrameStrobe_O(Tile_X4Y5_FrameStrobe_O)
	);


	LUT4AB Tile_X6Y5_LUT4AB (
	.N1END(Tile_X6Y6_N1BEG[3:0]),
	.N2MID(Tile_X6Y6_N2BEG[7:0]),
	.N2END(Tile_X6Y6_N2BEGb[7:0]),
	.N4END(Tile_X6Y6_N4BEG[15:0]),
	.NN4END(Tile_X6Y6_NN4BEG[15:0]),
	.Ci(Tile_X6Y6_Co[0:0]),
	.E1END(Tile_X5Y5_E1BEG[3:0]),
	.E2MID(Tile_X5Y5_E2BEG[7:0]),
	.E2END(Tile_X5Y5_E2BEGb[7:0]),
	.EE4END(Tile_X5Y5_EE4BEG[15:0]),
	.E6END(Tile_X5Y5_E6BEG[11:0]),
	.S1END(Tile_X6Y4_S1BEG[3:0]),
	.S2MID(Tile_X6Y4_S2BEG[7:0]),
	.S2END(Tile_X6Y4_S2BEGb[7:0]),
	.S4END(Tile_X6Y4_S4BEG[15:0]),
	.SS4END(Tile_X6Y4_SS4BEG[15:0]),
	.W1END(Tile_X7Y5_W1BEG[3:0]),
	.W2MID(Tile_X7Y5_W2BEG[7:0]),
	.W2END(Tile_X7Y5_W2BEGb[7:0]),
	.WW4END(Tile_X7Y5_WW4BEG[15:0]),
	.W6END(Tile_X7Y5_W6BEG[11:0]),
	.N1BEG(Tile_X6Y5_N1BEG[3:0]),
	.N2BEG(Tile_X6Y5_N2BEG[7:0]),
	.N2BEGb(Tile_X6Y5_N2BEGb[7:0]),
	.N4BEG(Tile_X6Y5_N4BEG[15:0]),
	.NN4BEG(Tile_X6Y5_NN4BEG[15:0]),
	.Co(Tile_X6Y5_Co[0:0]),
	.E1BEG(Tile_X6Y5_E1BEG[3:0]),
	.E2BEG(Tile_X6Y5_E2BEG[7:0]),
	.E2BEGb(Tile_X6Y5_E2BEGb[7:0]),
	.EE4BEG(Tile_X6Y5_EE4BEG[15:0]),
	.E6BEG(Tile_X6Y5_E6BEG[11:0]),
	.S1BEG(Tile_X6Y5_S1BEG[3:0]),
	.S2BEG(Tile_X6Y5_S2BEG[7:0]),
	.S2BEGb(Tile_X6Y5_S2BEGb[7:0]),
	.S4BEG(Tile_X6Y5_S4BEG[15:0]),
	.SS4BEG(Tile_X6Y5_SS4BEG[15:0]),
	.W1BEG(Tile_X6Y5_W1BEG[3:0]),
	.W2BEG(Tile_X6Y5_W2BEG[7:0]),
	.W2BEGb(Tile_X6Y5_W2BEGb[7:0]),
	.WW4BEG(Tile_X6Y5_WW4BEG[15:0]),
	.W6BEG(Tile_X6Y5_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X6Y6_UserCLKo),
	.UserCLKo(Tile_X6Y5_UserCLKo),
	.FrameData(Tile_X5Y5_FrameData_O), 
	.FrameData_O(Tile_X6Y5_FrameData_O), 
	.FrameStrobe(Tile_X6Y6_FrameStrobe_O),
	.FrameStrobe_O(Tile_X6Y5_FrameStrobe_O)
	);

	LUT4AB Tile_X7Y5_LUT4AB (
	.N1END(Tile_X7Y6_N1BEG[3:0]),
	.N2MID(Tile_X7Y6_N2BEG[7:0]),
	.N2END(Tile_X7Y6_N2BEGb[7:0]),
	.N4END(Tile_X7Y6_N4BEG[15:0]),
	.NN4END(Tile_X7Y6_NN4BEG[15:0]),
	.Ci(Tile_X7Y6_Co[0:0]),
	.E1END(Tile_X6Y5_E1BEG[3:0]),
	.E2MID(Tile_X6Y5_E2BEG[7:0]),
	.E2END(Tile_X6Y5_E2BEGb[7:0]),
	.EE4END(Tile_X6Y5_EE4BEG[15:0]),
	.E6END(Tile_X6Y5_E6BEG[11:0]),
	.S1END(Tile_X7Y4_S1BEG[3:0]),
	.S2MID(Tile_X7Y4_S2BEG[7:0]),
	.S2END(Tile_X7Y4_S2BEGb[7:0]),
	.S4END(Tile_X7Y4_S4BEG[15:0]),
	.SS4END(Tile_X7Y4_SS4BEG[15:0]),
	.W1END(Tile_X8Y5_W1BEG[3:0]),
	.W2MID(Tile_X8Y5_W2BEG[7:0]),
	.W2END(Tile_X8Y5_W2BEGb[7:0]),
	.WW4END(Tile_X8Y5_WW4BEG[15:0]),
	.W6END(Tile_X8Y5_W6BEG[11:0]),
	.N1BEG(Tile_X7Y5_N1BEG[3:0]),
	.N2BEG(Tile_X7Y5_N2BEG[7:0]),
	.N2BEGb(Tile_X7Y5_N2BEGb[7:0]),
	.N4BEG(Tile_X7Y5_N4BEG[15:0]),
	.NN4BEG(Tile_X7Y5_NN4BEG[15:0]),
	.Co(Tile_X7Y5_Co[0:0]),
	.E1BEG(Tile_X7Y5_E1BEG[3:0]),
	.E2BEG(Tile_X7Y5_E2BEG[7:0]),
	.E2BEGb(Tile_X7Y5_E2BEGb[7:0]),
	.EE4BEG(Tile_X7Y5_EE4BEG[15:0]),
	.E6BEG(Tile_X7Y5_E6BEG[11:0]),
	.S1BEG(Tile_X7Y5_S1BEG[3:0]),
	.S2BEG(Tile_X7Y5_S2BEG[7:0]),
	.S2BEGb(Tile_X7Y5_S2BEGb[7:0]),
	.S4BEG(Tile_X7Y5_S4BEG[15:0]),
	.SS4BEG(Tile_X7Y5_SS4BEG[15:0]),
	.W1BEG(Tile_X7Y5_W1BEG[3:0]),
	.W2BEG(Tile_X7Y5_W2BEG[7:0]),
	.W2BEGb(Tile_X7Y5_W2BEGb[7:0]),
	.WW4BEG(Tile_X7Y5_WW4BEG[15:0]),
	.W6BEG(Tile_X7Y5_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X7Y6_UserCLKo),
	.UserCLKo(Tile_X7Y5_UserCLKo),
	.FrameData(Tile_X6Y5_FrameData_O), 
	.FrameData_O(Tile_X7Y5_FrameData_O), 
	.FrameStrobe(Tile_X7Y6_FrameStrobe_O),
	.FrameStrobe_O(Tile_X7Y5_FrameStrobe_O)
	);

	LUT4AB Tile_X8Y5_LUT4AB (
	.N1END(Tile_X8Y6_N1BEG[3:0]),
	.N2MID(Tile_X8Y6_N2BEG[7:0]),
	.N2END(Tile_X8Y6_N2BEGb[7:0]),
	.N4END(Tile_X8Y6_N4BEG[15:0]),
	.NN4END(Tile_X8Y6_NN4BEG[15:0]),
	.Ci(Tile_X8Y6_Co[0:0]),
	.E1END(Tile_X7Y5_E1BEG[3:0]),
	.E2MID(Tile_X7Y5_E2BEG[7:0]),
	.E2END(Tile_X7Y5_E2BEGb[7:0]),
	.EE4END(Tile_X7Y5_EE4BEG[15:0]),
	.E6END(Tile_X7Y5_E6BEG[11:0]),
	.S1END(Tile_X8Y4_S1BEG[3:0]),
	.S2MID(Tile_X8Y4_S2BEG[7:0]),
	.S2END(Tile_X8Y4_S2BEGb[7:0]),
	.S4END(Tile_X8Y4_S4BEG[15:0]),
	.SS4END(Tile_X8Y4_SS4BEG[15:0]),
	.W1END(Tile_X9Y5_W1BEG[3:0]),
	.W2MID(Tile_X9Y5_W2BEG[7:0]),
	.W2END(Tile_X9Y5_W2BEGb[7:0]),
	.WW4END(Tile_X9Y5_WW4BEG[15:0]),
	.W6END(Tile_X9Y5_W6BEG[11:0]),
	.N1BEG(Tile_X8Y5_N1BEG[3:0]),
	.N2BEG(Tile_X8Y5_N2BEG[7:0]),
	.N2BEGb(Tile_X8Y5_N2BEGb[7:0]),
	.N4BEG(Tile_X8Y5_N4BEG[15:0]),
	.NN4BEG(Tile_X8Y5_NN4BEG[15:0]),
	.Co(Tile_X8Y5_Co[0:0]),
	.E1BEG(Tile_X8Y5_E1BEG[3:0]),
	.E2BEG(Tile_X8Y5_E2BEG[7:0]),
	.E2BEGb(Tile_X8Y5_E2BEGb[7:0]),
	.EE4BEG(Tile_X8Y5_EE4BEG[15:0]),
	.E6BEG(Tile_X8Y5_E6BEG[11:0]),
	.S1BEG(Tile_X8Y5_S1BEG[3:0]),
	.S2BEG(Tile_X8Y5_S2BEG[7:0]),
	.S2BEGb(Tile_X8Y5_S2BEGb[7:0]),
	.S4BEG(Tile_X8Y5_S4BEG[15:0]),
	.SS4BEG(Tile_X8Y5_SS4BEG[15:0]),
	.W1BEG(Tile_X8Y5_W1BEG[3:0]),
	.W2BEG(Tile_X8Y5_W2BEG[7:0]),
	.W2BEGb(Tile_X8Y5_W2BEGb[7:0]),
	.WW4BEG(Tile_X8Y5_WW4BEG[15:0]),
	.W6BEG(Tile_X8Y5_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X8Y6_UserCLKo),
	.UserCLKo(Tile_X8Y5_UserCLKo),
	.FrameData(Tile_X7Y5_FrameData_O), 
	.FrameData_O(Tile_X8Y5_FrameData_O), 
	.FrameStrobe(Tile_X8Y6_FrameStrobe_O),
	.FrameStrobe_O(Tile_X8Y5_FrameStrobe_O)
	);


	LUT4AB Tile_X10Y5_LUT4AB (
	.N1END(Tile_X10Y6_N1BEG[3:0]),
	.N2MID(Tile_X10Y6_N2BEG[7:0]),
	.N2END(Tile_X10Y6_N2BEGb[7:0]),
	.N4END(Tile_X10Y6_N4BEG[15:0]),
	.NN4END(Tile_X10Y6_NN4BEG[15:0]),
	.Ci(Tile_X10Y6_Co[0:0]),
	.E1END(Tile_X9Y5_E1BEG[3:0]),
	.E2MID(Tile_X9Y5_E2BEG[7:0]),
	.E2END(Tile_X9Y5_E2BEGb[7:0]),
	.EE4END(Tile_X9Y5_EE4BEG[15:0]),
	.E6END(Tile_X9Y5_E6BEG[11:0]),
	.S1END(Tile_X10Y4_S1BEG[3:0]),
	.S2MID(Tile_X10Y4_S2BEG[7:0]),
	.S2END(Tile_X10Y4_S2BEGb[7:0]),
	.S4END(Tile_X10Y4_S4BEG[15:0]),
	.SS4END(Tile_X10Y4_SS4BEG[15:0]),
	.W1END(Tile_X11Y5_W1BEG[3:0]),
	.W2MID(Tile_X11Y5_W2BEG[7:0]),
	.W2END(Tile_X11Y5_W2BEGb[7:0]),
	.WW4END(Tile_X11Y5_WW4BEG[15:0]),
	.W6END(Tile_X11Y5_W6BEG[11:0]),
	.N1BEG(Tile_X10Y5_N1BEG[3:0]),
	.N2BEG(Tile_X10Y5_N2BEG[7:0]),
	.N2BEGb(Tile_X10Y5_N2BEGb[7:0]),
	.N4BEG(Tile_X10Y5_N4BEG[15:0]),
	.NN4BEG(Tile_X10Y5_NN4BEG[15:0]),
	.Co(Tile_X10Y5_Co[0:0]),
	.E1BEG(Tile_X10Y5_E1BEG[3:0]),
	.E2BEG(Tile_X10Y5_E2BEG[7:0]),
	.E2BEGb(Tile_X10Y5_E2BEGb[7:0]),
	.EE4BEG(Tile_X10Y5_EE4BEG[15:0]),
	.E6BEG(Tile_X10Y5_E6BEG[11:0]),
	.S1BEG(Tile_X10Y5_S1BEG[3:0]),
	.S2BEG(Tile_X10Y5_S2BEG[7:0]),
	.S2BEGb(Tile_X10Y5_S2BEGb[7:0]),
	.S4BEG(Tile_X10Y5_S4BEG[15:0]),
	.SS4BEG(Tile_X10Y5_SS4BEG[15:0]),
	.W1BEG(Tile_X10Y5_W1BEG[3:0]),
	.W2BEG(Tile_X10Y5_W2BEG[7:0]),
	.W2BEGb(Tile_X10Y5_W2BEGb[7:0]),
	.WW4BEG(Tile_X10Y5_WW4BEG[15:0]),
	.W6BEG(Tile_X10Y5_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X10Y6_UserCLKo),
	.UserCLKo(Tile_X10Y5_UserCLKo),
	.FrameData(Tile_X9Y5_FrameData_O), 
	.FrameData_O(Tile_X10Y5_FrameData_O), 
	.FrameStrobe(Tile_X10Y6_FrameStrobe_O),
	.FrameStrobe_O(Tile_X10Y5_FrameStrobe_O)
	);

	E_CPU_IO Tile_X11Y5_E_CPU_IO (
	.E1END(Tile_X10Y5_E1BEG[3:0]),
	.E2MID(Tile_X10Y5_E2BEG[7:0]),
	.E2END(Tile_X10Y5_E2BEGb[7:0]),
	.EE4END(Tile_X10Y5_EE4BEG[15:0]),
	.E6END(Tile_X10Y5_E6BEG[11:0]),
	.W1BEG(Tile_X11Y5_W1BEG[3:0]),
	.W2BEG(Tile_X11Y5_W2BEG[7:0]),
	.W2BEGb(Tile_X11Y5_W2BEGb[7:0]),
	.WW4BEG(Tile_X11Y5_WW4BEG[15:0]),
	.W6BEG(Tile_X11Y5_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X11Y5_OPA_I0),
	.OPA_I1(Tile_X11Y5_OPA_I1),
	.OPA_I2(Tile_X11Y5_OPA_I2),
	.OPA_I3(Tile_X11Y5_OPA_I3),
	.UserCLK(Tile_X11Y6_UserCLKo),
	.OPB_I0(Tile_X11Y5_OPB_I0),
	.OPB_I1(Tile_X11Y5_OPB_I1),
	.OPB_I2(Tile_X11Y5_OPB_I2),
	.OPB_I3(Tile_X11Y5_OPB_I3),
	.RES0_O0(Tile_X11Y5_RES0_O0),
	.RES0_O1(Tile_X11Y5_RES0_O1),
	.RES0_O2(Tile_X11Y5_RES0_O2),
	.RES0_O3(Tile_X11Y5_RES0_O3),
	.RES1_O0(Tile_X11Y5_RES1_O0),
	.RES1_O1(Tile_X11Y5_RES1_O1),
	.RES1_O2(Tile_X11Y5_RES1_O2),
	.RES1_O3(Tile_X11Y5_RES1_O3),
	.RES2_O0(Tile_X11Y5_RES2_O0),
	.RES2_O1(Tile_X11Y5_RES2_O1),
	.RES2_O2(Tile_X11Y5_RES2_O2),
	.RES2_O3(Tile_X11Y5_RES2_O3),
	.UserCLKo(Tile_X11Y5_UserCLKo),
	.FrameData(Tile_X10Y5_FrameData_O), 
	.FrameData_O(Tile_X11Y5_FrameData_O), 
	.FrameStrobe(Tile_X11Y6_FrameStrobe_O),
	.FrameStrobe_O(Tile_X11Y5_FrameStrobe_O)
	);

	W_CPU_IO Tile_X4Y6_W_CPU_IO (
	.W1END(Tile_X5Y6_W1BEG[3:0]),
	.W2MID(Tile_X5Y6_W2BEG[7:0]),
	.W2END(Tile_X5Y6_W2BEGb[7:0]),
	.WW4END(Tile_X5Y6_WW4BEG[15:0]),
	.W6END(Tile_X5Y6_W6BEG[11:0]),
	.E1BEG(Tile_X4Y6_E1BEG[3:0]),
	.E2BEG(Tile_X4Y6_E2BEG[7:0]),
	.E2BEGb(Tile_X4Y6_E2BEGb[7:0]),
	.EE4BEG(Tile_X4Y6_EE4BEG[15:0]),
	.E6BEG(Tile_X4Y6_E6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X4Y6_OPA_I0),
	.OPA_I1(Tile_X4Y6_OPA_I1),
	.OPA_I2(Tile_X4Y6_OPA_I2),
	.OPA_I3(Tile_X4Y6_OPA_I3),
	.UserCLK(Tile_X4Y7_UserCLKo),
	.OPB_I0(Tile_X4Y6_OPB_I0),
	.OPB_I1(Tile_X4Y6_OPB_I1),
	.OPB_I2(Tile_X4Y6_OPB_I2),
	.OPB_I3(Tile_X4Y6_OPB_I3),
	.RES0_O0(Tile_X4Y6_RES0_O0),
	.RES0_O1(Tile_X4Y6_RES0_O1),
	.RES0_O2(Tile_X4Y6_RES0_O2),
	.RES0_O3(Tile_X4Y6_RES0_O3),
	.RES1_O0(Tile_X4Y6_RES1_O0),
	.RES1_O1(Tile_X4Y6_RES1_O1),
	.RES1_O2(Tile_X4Y6_RES1_O2),
	.RES1_O3(Tile_X4Y6_RES1_O3),
	.RES2_O0(Tile_X4Y6_RES2_O0),
	.RES2_O1(Tile_X4Y6_RES2_O1),
	.RES2_O2(Tile_X4Y6_RES2_O2),
	.RES2_O3(Tile_X4Y6_RES2_O3),
	.UserCLKo(Tile_X4Y6_UserCLKo),
	.FrameData(Tile_Y6_FrameData), 
	.FrameData_O(Tile_X4Y6_FrameData_O), 
	.FrameStrobe(Tile_X4Y7_FrameStrobe_O),
	.FrameStrobe_O(Tile_X4Y6_FrameStrobe_O)
	);


	LUT4AB Tile_X6Y6_LUT4AB (
	.N1END(Tile_X6Y7_N1BEG[3:0]),
	.N2MID(Tile_X6Y7_N2BEG[7:0]),
	.N2END(Tile_X6Y7_N2BEGb[7:0]),
	.N4END(Tile_X6Y7_N4BEG[15:0]),
	.NN4END(Tile_X6Y7_NN4BEG[15:0]),
	.Ci(Tile_X6Y7_Co[0:0]),
	.E1END(Tile_X5Y6_E1BEG[3:0]),
	.E2MID(Tile_X5Y6_E2BEG[7:0]),
	.E2END(Tile_X5Y6_E2BEGb[7:0]),
	.EE4END(Tile_X5Y6_EE4BEG[15:0]),
	.E6END(Tile_X5Y6_E6BEG[11:0]),
	.S1END(Tile_X6Y5_S1BEG[3:0]),
	.S2MID(Tile_X6Y5_S2BEG[7:0]),
	.S2END(Tile_X6Y5_S2BEGb[7:0]),
	.S4END(Tile_X6Y5_S4BEG[15:0]),
	.SS4END(Tile_X6Y5_SS4BEG[15:0]),
	.W1END(Tile_X7Y6_W1BEG[3:0]),
	.W2MID(Tile_X7Y6_W2BEG[7:0]),
	.W2END(Tile_X7Y6_W2BEGb[7:0]),
	.WW4END(Tile_X7Y6_WW4BEG[15:0]),
	.W6END(Tile_X7Y6_W6BEG[11:0]),
	.N1BEG(Tile_X6Y6_N1BEG[3:0]),
	.N2BEG(Tile_X6Y6_N2BEG[7:0]),
	.N2BEGb(Tile_X6Y6_N2BEGb[7:0]),
	.N4BEG(Tile_X6Y6_N4BEG[15:0]),
	.NN4BEG(Tile_X6Y6_NN4BEG[15:0]),
	.Co(Tile_X6Y6_Co[0:0]),
	.E1BEG(Tile_X6Y6_E1BEG[3:0]),
	.E2BEG(Tile_X6Y6_E2BEG[7:0]),
	.E2BEGb(Tile_X6Y6_E2BEGb[7:0]),
	.EE4BEG(Tile_X6Y6_EE4BEG[15:0]),
	.E6BEG(Tile_X6Y6_E6BEG[11:0]),
	.S1BEG(Tile_X6Y6_S1BEG[3:0]),
	.S2BEG(Tile_X6Y6_S2BEG[7:0]),
	.S2BEGb(Tile_X6Y6_S2BEGb[7:0]),
	.S4BEG(Tile_X6Y6_S4BEG[15:0]),
	.SS4BEG(Tile_X6Y6_SS4BEG[15:0]),
	.W1BEG(Tile_X6Y6_W1BEG[3:0]),
	.W2BEG(Tile_X6Y6_W2BEG[7:0]),
	.W2BEGb(Tile_X6Y6_W2BEGb[7:0]),
	.WW4BEG(Tile_X6Y6_WW4BEG[15:0]),
	.W6BEG(Tile_X6Y6_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X6Y7_UserCLKo),
	.UserCLKo(Tile_X6Y6_UserCLKo),
	.FrameData(Tile_X5Y6_FrameData_O), 
	.FrameData_O(Tile_X6Y6_FrameData_O), 
	.FrameStrobe(Tile_X6Y7_FrameStrobe_O),
	.FrameStrobe_O(Tile_X6Y6_FrameStrobe_O)
	);

	LUT4AB Tile_X7Y6_LUT4AB (
	.N1END(Tile_X7Y7_N1BEG[3:0]),
	.N2MID(Tile_X7Y7_N2BEG[7:0]),
	.N2END(Tile_X7Y7_N2BEGb[7:0]),
	.N4END(Tile_X7Y7_N4BEG[15:0]),
	.NN4END(Tile_X7Y7_NN4BEG[15:0]),
	.Ci(Tile_X7Y7_Co[0:0]),
	.E1END(Tile_X6Y6_E1BEG[3:0]),
	.E2MID(Tile_X6Y6_E2BEG[7:0]),
	.E2END(Tile_X6Y6_E2BEGb[7:0]),
	.EE4END(Tile_X6Y6_EE4BEG[15:0]),
	.E6END(Tile_X6Y6_E6BEG[11:0]),
	.S1END(Tile_X7Y5_S1BEG[3:0]),
	.S2MID(Tile_X7Y5_S2BEG[7:0]),
	.S2END(Tile_X7Y5_S2BEGb[7:0]),
	.S4END(Tile_X7Y5_S4BEG[15:0]),
	.SS4END(Tile_X7Y5_SS4BEG[15:0]),
	.W1END(Tile_X8Y6_W1BEG[3:0]),
	.W2MID(Tile_X8Y6_W2BEG[7:0]),
	.W2END(Tile_X8Y6_W2BEGb[7:0]),
	.WW4END(Tile_X8Y6_WW4BEG[15:0]),
	.W6END(Tile_X8Y6_W6BEG[11:0]),
	.N1BEG(Tile_X7Y6_N1BEG[3:0]),
	.N2BEG(Tile_X7Y6_N2BEG[7:0]),
	.N2BEGb(Tile_X7Y6_N2BEGb[7:0]),
	.N4BEG(Tile_X7Y6_N4BEG[15:0]),
	.NN4BEG(Tile_X7Y6_NN4BEG[15:0]),
	.Co(Tile_X7Y6_Co[0:0]),
	.E1BEG(Tile_X7Y6_E1BEG[3:0]),
	.E2BEG(Tile_X7Y6_E2BEG[7:0]),
	.E2BEGb(Tile_X7Y6_E2BEGb[7:0]),
	.EE4BEG(Tile_X7Y6_EE4BEG[15:0]),
	.E6BEG(Tile_X7Y6_E6BEG[11:0]),
	.S1BEG(Tile_X7Y6_S1BEG[3:0]),
	.S2BEG(Tile_X7Y6_S2BEG[7:0]),
	.S2BEGb(Tile_X7Y6_S2BEGb[7:0]),
	.S4BEG(Tile_X7Y6_S4BEG[15:0]),
	.SS4BEG(Tile_X7Y6_SS4BEG[15:0]),
	.W1BEG(Tile_X7Y6_W1BEG[3:0]),
	.W2BEG(Tile_X7Y6_W2BEG[7:0]),
	.W2BEGb(Tile_X7Y6_W2BEGb[7:0]),
	.WW4BEG(Tile_X7Y6_WW4BEG[15:0]),
	.W6BEG(Tile_X7Y6_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X7Y7_UserCLKo),
	.UserCLKo(Tile_X7Y6_UserCLKo),
	.FrameData(Tile_X6Y6_FrameData_O), 
	.FrameData_O(Tile_X7Y6_FrameData_O), 
	.FrameStrobe(Tile_X7Y7_FrameStrobe_O),
	.FrameStrobe_O(Tile_X7Y6_FrameStrobe_O)
	);

	LUT4AB Tile_X8Y6_LUT4AB (
	.N1END(Tile_X8Y7_N1BEG[3:0]),
	.N2MID(Tile_X8Y7_N2BEG[7:0]),
	.N2END(Tile_X8Y7_N2BEGb[7:0]),
	.N4END(Tile_X8Y7_N4BEG[15:0]),
	.NN4END(Tile_X8Y7_NN4BEG[15:0]),
	.Ci(Tile_X8Y7_Co[0:0]),
	.E1END(Tile_X7Y6_E1BEG[3:0]),
	.E2MID(Tile_X7Y6_E2BEG[7:0]),
	.E2END(Tile_X7Y6_E2BEGb[7:0]),
	.EE4END(Tile_X7Y6_EE4BEG[15:0]),
	.E6END(Tile_X7Y6_E6BEG[11:0]),
	.S1END(Tile_X8Y5_S1BEG[3:0]),
	.S2MID(Tile_X8Y5_S2BEG[7:0]),
	.S2END(Tile_X8Y5_S2BEGb[7:0]),
	.S4END(Tile_X8Y5_S4BEG[15:0]),
	.SS4END(Tile_X8Y5_SS4BEG[15:0]),
	.W1END(Tile_X9Y6_W1BEG[3:0]),
	.W2MID(Tile_X9Y6_W2BEG[7:0]),
	.W2END(Tile_X9Y6_W2BEGb[7:0]),
	.WW4END(Tile_X9Y6_WW4BEG[15:0]),
	.W6END(Tile_X9Y6_W6BEG[11:0]),
	.N1BEG(Tile_X8Y6_N1BEG[3:0]),
	.N2BEG(Tile_X8Y6_N2BEG[7:0]),
	.N2BEGb(Tile_X8Y6_N2BEGb[7:0]),
	.N4BEG(Tile_X8Y6_N4BEG[15:0]),
	.NN4BEG(Tile_X8Y6_NN4BEG[15:0]),
	.Co(Tile_X8Y6_Co[0:0]),
	.E1BEG(Tile_X8Y6_E1BEG[3:0]),
	.E2BEG(Tile_X8Y6_E2BEG[7:0]),
	.E2BEGb(Tile_X8Y6_E2BEGb[7:0]),
	.EE4BEG(Tile_X8Y6_EE4BEG[15:0]),
	.E6BEG(Tile_X8Y6_E6BEG[11:0]),
	.S1BEG(Tile_X8Y6_S1BEG[3:0]),
	.S2BEG(Tile_X8Y6_S2BEG[7:0]),
	.S2BEGb(Tile_X8Y6_S2BEGb[7:0]),
	.S4BEG(Tile_X8Y6_S4BEG[15:0]),
	.SS4BEG(Tile_X8Y6_SS4BEG[15:0]),
	.W1BEG(Tile_X8Y6_W1BEG[3:0]),
	.W2BEG(Tile_X8Y6_W2BEG[7:0]),
	.W2BEGb(Tile_X8Y6_W2BEGb[7:0]),
	.WW4BEG(Tile_X8Y6_WW4BEG[15:0]),
	.W6BEG(Tile_X8Y6_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X8Y7_UserCLKo),
	.UserCLKo(Tile_X8Y6_UserCLKo),
	.FrameData(Tile_X7Y6_FrameData_O), 
	.FrameData_O(Tile_X8Y6_FrameData_O), 
	.FrameStrobe(Tile_X8Y7_FrameStrobe_O),
	.FrameStrobe_O(Tile_X8Y6_FrameStrobe_O)
	);


	LUT4AB Tile_X10Y6_LUT4AB (
	.N1END(Tile_X10Y7_N1BEG[3:0]),
	.N2MID(Tile_X10Y7_N2BEG[7:0]),
	.N2END(Tile_X10Y7_N2BEGb[7:0]),
	.N4END(Tile_X10Y7_N4BEG[15:0]),
	.NN4END(Tile_X10Y7_NN4BEG[15:0]),
	.Ci(Tile_X10Y7_Co[0:0]),
	.E1END(Tile_X9Y6_E1BEG[3:0]),
	.E2MID(Tile_X9Y6_E2BEG[7:0]),
	.E2END(Tile_X9Y6_E2BEGb[7:0]),
	.EE4END(Tile_X9Y6_EE4BEG[15:0]),
	.E6END(Tile_X9Y6_E6BEG[11:0]),
	.S1END(Tile_X10Y5_S1BEG[3:0]),
	.S2MID(Tile_X10Y5_S2BEG[7:0]),
	.S2END(Tile_X10Y5_S2BEGb[7:0]),
	.S4END(Tile_X10Y5_S4BEG[15:0]),
	.SS4END(Tile_X10Y5_SS4BEG[15:0]),
	.W1END(Tile_X11Y6_W1BEG[3:0]),
	.W2MID(Tile_X11Y6_W2BEG[7:0]),
	.W2END(Tile_X11Y6_W2BEGb[7:0]),
	.WW4END(Tile_X11Y6_WW4BEG[15:0]),
	.W6END(Tile_X11Y6_W6BEG[11:0]),
	.N1BEG(Tile_X10Y6_N1BEG[3:0]),
	.N2BEG(Tile_X10Y6_N2BEG[7:0]),
	.N2BEGb(Tile_X10Y6_N2BEGb[7:0]),
	.N4BEG(Tile_X10Y6_N4BEG[15:0]),
	.NN4BEG(Tile_X10Y6_NN4BEG[15:0]),
	.Co(Tile_X10Y6_Co[0:0]),
	.E1BEG(Tile_X10Y6_E1BEG[3:0]),
	.E2BEG(Tile_X10Y6_E2BEG[7:0]),
	.E2BEGb(Tile_X10Y6_E2BEGb[7:0]),
	.EE4BEG(Tile_X10Y6_EE4BEG[15:0]),
	.E6BEG(Tile_X10Y6_E6BEG[11:0]),
	.S1BEG(Tile_X10Y6_S1BEG[3:0]),
	.S2BEG(Tile_X10Y6_S2BEG[7:0]),
	.S2BEGb(Tile_X10Y6_S2BEGb[7:0]),
	.S4BEG(Tile_X10Y6_S4BEG[15:0]),
	.SS4BEG(Tile_X10Y6_SS4BEG[15:0]),
	.W1BEG(Tile_X10Y6_W1BEG[3:0]),
	.W2BEG(Tile_X10Y6_W2BEG[7:0]),
	.W2BEGb(Tile_X10Y6_W2BEGb[7:0]),
	.WW4BEG(Tile_X10Y6_WW4BEG[15:0]),
	.W6BEG(Tile_X10Y6_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X10Y7_UserCLKo),
	.UserCLKo(Tile_X10Y6_UserCLKo),
	.FrameData(Tile_X9Y6_FrameData_O), 
	.FrameData_O(Tile_X10Y6_FrameData_O), 
	.FrameStrobe(Tile_X10Y7_FrameStrobe_O),
	.FrameStrobe_O(Tile_X10Y6_FrameStrobe_O)
	);

	E_CPU_IO Tile_X11Y6_E_CPU_IO (
	.E1END(Tile_X10Y6_E1BEG[3:0]),
	.E2MID(Tile_X10Y6_E2BEG[7:0]),
	.E2END(Tile_X10Y6_E2BEGb[7:0]),
	.EE4END(Tile_X10Y6_EE4BEG[15:0]),
	.E6END(Tile_X10Y6_E6BEG[11:0]),
	.W1BEG(Tile_X11Y6_W1BEG[3:0]),
	.W2BEG(Tile_X11Y6_W2BEG[7:0]),
	.W2BEGb(Tile_X11Y6_W2BEGb[7:0]),
	.WW4BEG(Tile_X11Y6_WW4BEG[15:0]),
	.W6BEG(Tile_X11Y6_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X11Y6_OPA_I0),
	.OPA_I1(Tile_X11Y6_OPA_I1),
	.OPA_I2(Tile_X11Y6_OPA_I2),
	.OPA_I3(Tile_X11Y6_OPA_I3),
	.UserCLK(Tile_X11Y7_UserCLKo),
	.OPB_I0(Tile_X11Y6_OPB_I0),
	.OPB_I1(Tile_X11Y6_OPB_I1),
	.OPB_I2(Tile_X11Y6_OPB_I2),
	.OPB_I3(Tile_X11Y6_OPB_I3),
	.RES0_O0(Tile_X11Y6_RES0_O0),
	.RES0_O1(Tile_X11Y6_RES0_O1),
	.RES0_O2(Tile_X11Y6_RES0_O2),
	.RES0_O3(Tile_X11Y6_RES0_O3),
	.RES1_O0(Tile_X11Y6_RES1_O0),
	.RES1_O1(Tile_X11Y6_RES1_O1),
	.RES1_O2(Tile_X11Y6_RES1_O2),
	.RES1_O3(Tile_X11Y6_RES1_O3),
	.RES2_O0(Tile_X11Y6_RES2_O0),
	.RES2_O1(Tile_X11Y6_RES2_O1),
	.RES2_O2(Tile_X11Y6_RES2_O2),
	.RES2_O3(Tile_X11Y6_RES2_O3),
	.UserCLKo(Tile_X11Y6_UserCLKo),
	.FrameData(Tile_X10Y6_FrameData_O), 
	.FrameData_O(Tile_X11Y6_FrameData_O), 
	.FrameStrobe(Tile_X11Y7_FrameStrobe_O),
	.FrameStrobe_O(Tile_X11Y6_FrameStrobe_O)
	);

	W_CPU_IO Tile_X4Y7_W_CPU_IO (
	.W1END(Tile_X5Y7_W1BEG[3:0]),
	.W2MID(Tile_X5Y7_W2BEG[7:0]),
	.W2END(Tile_X5Y7_W2BEGb[7:0]),
	.WW4END(Tile_X5Y7_WW4BEG[15:0]),
	.W6END(Tile_X5Y7_W6BEG[11:0]),
	.E1BEG(Tile_X4Y7_E1BEG[3:0]),
	.E2BEG(Tile_X4Y7_E2BEG[7:0]),
	.E2BEGb(Tile_X4Y7_E2BEGb[7:0]),
	.EE4BEG(Tile_X4Y7_EE4BEG[15:0]),
	.E6BEG(Tile_X4Y7_E6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X4Y7_OPA_I0),
	.OPA_I1(Tile_X4Y7_OPA_I1),
	.OPA_I2(Tile_X4Y7_OPA_I2),
	.OPA_I3(Tile_X4Y7_OPA_I3),
	.UserCLK(Tile_X4Y8_UserCLKo),
	.OPB_I0(Tile_X4Y7_OPB_I0),
	.OPB_I1(Tile_X4Y7_OPB_I1),
	.OPB_I2(Tile_X4Y7_OPB_I2),
	.OPB_I3(Tile_X4Y7_OPB_I3),
	.RES0_O0(Tile_X4Y7_RES0_O0),
	.RES0_O1(Tile_X4Y7_RES0_O1),
	.RES0_O2(Tile_X4Y7_RES0_O2),
	.RES0_O3(Tile_X4Y7_RES0_O3),
	.RES1_O0(Tile_X4Y7_RES1_O0),
	.RES1_O1(Tile_X4Y7_RES1_O1),
	.RES1_O2(Tile_X4Y7_RES1_O2),
	.RES1_O3(Tile_X4Y7_RES1_O3),
	.RES2_O0(Tile_X4Y7_RES2_O0),
	.RES2_O1(Tile_X4Y7_RES2_O1),
	.RES2_O2(Tile_X4Y7_RES2_O2),
	.RES2_O3(Tile_X4Y7_RES2_O3),
	.UserCLKo(Tile_X4Y7_UserCLKo),
	.FrameData(Tile_Y7_FrameData), 
	.FrameData_O(Tile_X4Y7_FrameData_O), 
	.FrameStrobe(Tile_X4Y8_FrameStrobe_O),
	.FrameStrobe_O(Tile_X4Y7_FrameStrobe_O)
	);


	LUT4AB Tile_X6Y7_LUT4AB (
	.N1END(Tile_X6Y8_N1BEG[3:0]),
	.N2MID(Tile_X6Y8_N2BEG[7:0]),
	.N2END(Tile_X6Y8_N2BEGb[7:0]),
	.N4END(Tile_X6Y8_N4BEG[15:0]),
	.NN4END(Tile_X6Y8_NN4BEG[15:0]),
	.Ci(Tile_X6Y8_Co[0:0]),
	.E1END(Tile_X5Y7_E1BEG[3:0]),
	.E2MID(Tile_X5Y7_E2BEG[7:0]),
	.E2END(Tile_X5Y7_E2BEGb[7:0]),
	.EE4END(Tile_X5Y7_EE4BEG[15:0]),
	.E6END(Tile_X5Y7_E6BEG[11:0]),
	.S1END(Tile_X6Y6_S1BEG[3:0]),
	.S2MID(Tile_X6Y6_S2BEG[7:0]),
	.S2END(Tile_X6Y6_S2BEGb[7:0]),
	.S4END(Tile_X6Y6_S4BEG[15:0]),
	.SS4END(Tile_X6Y6_SS4BEG[15:0]),
	.W1END(Tile_X7Y7_W1BEG[3:0]),
	.W2MID(Tile_X7Y7_W2BEG[7:0]),
	.W2END(Tile_X7Y7_W2BEGb[7:0]),
	.WW4END(Tile_X7Y7_WW4BEG[15:0]),
	.W6END(Tile_X7Y7_W6BEG[11:0]),
	.N1BEG(Tile_X6Y7_N1BEG[3:0]),
	.N2BEG(Tile_X6Y7_N2BEG[7:0]),
	.N2BEGb(Tile_X6Y7_N2BEGb[7:0]),
	.N4BEG(Tile_X6Y7_N4BEG[15:0]),
	.NN4BEG(Tile_X6Y7_NN4BEG[15:0]),
	.Co(Tile_X6Y7_Co[0:0]),
	.E1BEG(Tile_X6Y7_E1BEG[3:0]),
	.E2BEG(Tile_X6Y7_E2BEG[7:0]),
	.E2BEGb(Tile_X6Y7_E2BEGb[7:0]),
	.EE4BEG(Tile_X6Y7_EE4BEG[15:0]),
	.E6BEG(Tile_X6Y7_E6BEG[11:0]),
	.S1BEG(Tile_X6Y7_S1BEG[3:0]),
	.S2BEG(Tile_X6Y7_S2BEG[7:0]),
	.S2BEGb(Tile_X6Y7_S2BEGb[7:0]),
	.S4BEG(Tile_X6Y7_S4BEG[15:0]),
	.SS4BEG(Tile_X6Y7_SS4BEG[15:0]),
	.W1BEG(Tile_X6Y7_W1BEG[3:0]),
	.W2BEG(Tile_X6Y7_W2BEG[7:0]),
	.W2BEGb(Tile_X6Y7_W2BEGb[7:0]),
	.WW4BEG(Tile_X6Y7_WW4BEG[15:0]),
	.W6BEG(Tile_X6Y7_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X6Y8_UserCLKo),
	.UserCLKo(Tile_X6Y7_UserCLKo),
	.FrameData(Tile_X5Y7_FrameData_O), 
	.FrameData_O(Tile_X6Y7_FrameData_O), 
	.FrameStrobe(Tile_X6Y8_FrameStrobe_O),
	.FrameStrobe_O(Tile_X6Y7_FrameStrobe_O)
	);

	LUT4AB Tile_X7Y7_LUT4AB (
	.N1END(Tile_X7Y8_N1BEG[3:0]),
	.N2MID(Tile_X7Y8_N2BEG[7:0]),
	.N2END(Tile_X7Y8_N2BEGb[7:0]),
	.N4END(Tile_X7Y8_N4BEG[15:0]),
	.NN4END(Tile_X7Y8_NN4BEG[15:0]),
	.Ci(Tile_X7Y8_Co[0:0]),
	.E1END(Tile_X6Y7_E1BEG[3:0]),
	.E2MID(Tile_X6Y7_E2BEG[7:0]),
	.E2END(Tile_X6Y7_E2BEGb[7:0]),
	.EE4END(Tile_X6Y7_EE4BEG[15:0]),
	.E6END(Tile_X6Y7_E6BEG[11:0]),
	.S1END(Tile_X7Y6_S1BEG[3:0]),
	.S2MID(Tile_X7Y6_S2BEG[7:0]),
	.S2END(Tile_X7Y6_S2BEGb[7:0]),
	.S4END(Tile_X7Y6_S4BEG[15:0]),
	.SS4END(Tile_X7Y6_SS4BEG[15:0]),
	.W1END(Tile_X8Y7_W1BEG[3:0]),
	.W2MID(Tile_X8Y7_W2BEG[7:0]),
	.W2END(Tile_X8Y7_W2BEGb[7:0]),
	.WW4END(Tile_X8Y7_WW4BEG[15:0]),
	.W6END(Tile_X8Y7_W6BEG[11:0]),
	.N1BEG(Tile_X7Y7_N1BEG[3:0]),
	.N2BEG(Tile_X7Y7_N2BEG[7:0]),
	.N2BEGb(Tile_X7Y7_N2BEGb[7:0]),
	.N4BEG(Tile_X7Y7_N4BEG[15:0]),
	.NN4BEG(Tile_X7Y7_NN4BEG[15:0]),
	.Co(Tile_X7Y7_Co[0:0]),
	.E1BEG(Tile_X7Y7_E1BEG[3:0]),
	.E2BEG(Tile_X7Y7_E2BEG[7:0]),
	.E2BEGb(Tile_X7Y7_E2BEGb[7:0]),
	.EE4BEG(Tile_X7Y7_EE4BEG[15:0]),
	.E6BEG(Tile_X7Y7_E6BEG[11:0]),
	.S1BEG(Tile_X7Y7_S1BEG[3:0]),
	.S2BEG(Tile_X7Y7_S2BEG[7:0]),
	.S2BEGb(Tile_X7Y7_S2BEGb[7:0]),
	.S4BEG(Tile_X7Y7_S4BEG[15:0]),
	.SS4BEG(Tile_X7Y7_SS4BEG[15:0]),
	.W1BEG(Tile_X7Y7_W1BEG[3:0]),
	.W2BEG(Tile_X7Y7_W2BEG[7:0]),
	.W2BEGb(Tile_X7Y7_W2BEGb[7:0]),
	.WW4BEG(Tile_X7Y7_WW4BEG[15:0]),
	.W6BEG(Tile_X7Y7_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X7Y8_UserCLKo),
	.UserCLKo(Tile_X7Y7_UserCLKo),
	.FrameData(Tile_X6Y7_FrameData_O), 
	.FrameData_O(Tile_X7Y7_FrameData_O), 
	.FrameStrobe(Tile_X7Y8_FrameStrobe_O),
	.FrameStrobe_O(Tile_X7Y7_FrameStrobe_O)
	);

	LUT4AB Tile_X8Y7_LUT4AB (
	.N1END(Tile_X8Y8_N1BEG[3:0]),
	.N2MID(Tile_X8Y8_N2BEG[7:0]),
	.N2END(Tile_X8Y8_N2BEGb[7:0]),
	.N4END(Tile_X8Y8_N4BEG[15:0]),
	.NN4END(Tile_X8Y8_NN4BEG[15:0]),
	.Ci(Tile_X8Y8_Co[0:0]),
	.E1END(Tile_X7Y7_E1BEG[3:0]),
	.E2MID(Tile_X7Y7_E2BEG[7:0]),
	.E2END(Tile_X7Y7_E2BEGb[7:0]),
	.EE4END(Tile_X7Y7_EE4BEG[15:0]),
	.E6END(Tile_X7Y7_E6BEG[11:0]),
	.S1END(Tile_X8Y6_S1BEG[3:0]),
	.S2MID(Tile_X8Y6_S2BEG[7:0]),
	.S2END(Tile_X8Y6_S2BEGb[7:0]),
	.S4END(Tile_X8Y6_S4BEG[15:0]),
	.SS4END(Tile_X8Y6_SS4BEG[15:0]),
	.W1END(Tile_X9Y7_W1BEG[3:0]),
	.W2MID(Tile_X9Y7_W2BEG[7:0]),
	.W2END(Tile_X9Y7_W2BEGb[7:0]),
	.WW4END(Tile_X9Y7_WW4BEG[15:0]),
	.W6END(Tile_X9Y7_W6BEG[11:0]),
	.N1BEG(Tile_X8Y7_N1BEG[3:0]),
	.N2BEG(Tile_X8Y7_N2BEG[7:0]),
	.N2BEGb(Tile_X8Y7_N2BEGb[7:0]),
	.N4BEG(Tile_X8Y7_N4BEG[15:0]),
	.NN4BEG(Tile_X8Y7_NN4BEG[15:0]),
	.Co(Tile_X8Y7_Co[0:0]),
	.E1BEG(Tile_X8Y7_E1BEG[3:0]),
	.E2BEG(Tile_X8Y7_E2BEG[7:0]),
	.E2BEGb(Tile_X8Y7_E2BEGb[7:0]),
	.EE4BEG(Tile_X8Y7_EE4BEG[15:0]),
	.E6BEG(Tile_X8Y7_E6BEG[11:0]),
	.S1BEG(Tile_X8Y7_S1BEG[3:0]),
	.S2BEG(Tile_X8Y7_S2BEG[7:0]),
	.S2BEGb(Tile_X8Y7_S2BEGb[7:0]),
	.S4BEG(Tile_X8Y7_S4BEG[15:0]),
	.SS4BEG(Tile_X8Y7_SS4BEG[15:0]),
	.W1BEG(Tile_X8Y7_W1BEG[3:0]),
	.W2BEG(Tile_X8Y7_W2BEG[7:0]),
	.W2BEGb(Tile_X8Y7_W2BEGb[7:0]),
	.WW4BEG(Tile_X8Y7_WW4BEG[15:0]),
	.W6BEG(Tile_X8Y7_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X8Y8_UserCLKo),
	.UserCLKo(Tile_X8Y7_UserCLKo),
	.FrameData(Tile_X7Y7_FrameData_O), 
	.FrameData_O(Tile_X8Y7_FrameData_O), 
	.FrameStrobe(Tile_X8Y8_FrameStrobe_O),
	.FrameStrobe_O(Tile_X8Y7_FrameStrobe_O)
	);


	LUT4AB Tile_X10Y7_LUT4AB (
	.N1END(Tile_X10Y8_N1BEG[3:0]),
	.N2MID(Tile_X10Y8_N2BEG[7:0]),
	.N2END(Tile_X10Y8_N2BEGb[7:0]),
	.N4END(Tile_X10Y8_N4BEG[15:0]),
	.NN4END(Tile_X10Y8_NN4BEG[15:0]),
	.Ci(Tile_X10Y8_Co[0:0]),
	.E1END(Tile_X9Y7_E1BEG[3:0]),
	.E2MID(Tile_X9Y7_E2BEG[7:0]),
	.E2END(Tile_X9Y7_E2BEGb[7:0]),
	.EE4END(Tile_X9Y7_EE4BEG[15:0]),
	.E6END(Tile_X9Y7_E6BEG[11:0]),
	.S1END(Tile_X10Y6_S1BEG[3:0]),
	.S2MID(Tile_X10Y6_S2BEG[7:0]),
	.S2END(Tile_X10Y6_S2BEGb[7:0]),
	.S4END(Tile_X10Y6_S4BEG[15:0]),
	.SS4END(Tile_X10Y6_SS4BEG[15:0]),
	.W1END(Tile_X11Y7_W1BEG[3:0]),
	.W2MID(Tile_X11Y7_W2BEG[7:0]),
	.W2END(Tile_X11Y7_W2BEGb[7:0]),
	.WW4END(Tile_X11Y7_WW4BEG[15:0]),
	.W6END(Tile_X11Y7_W6BEG[11:0]),
	.N1BEG(Tile_X10Y7_N1BEG[3:0]),
	.N2BEG(Tile_X10Y7_N2BEG[7:0]),
	.N2BEGb(Tile_X10Y7_N2BEGb[7:0]),
	.N4BEG(Tile_X10Y7_N4BEG[15:0]),
	.NN4BEG(Tile_X10Y7_NN4BEG[15:0]),
	.Co(Tile_X10Y7_Co[0:0]),
	.E1BEG(Tile_X10Y7_E1BEG[3:0]),
	.E2BEG(Tile_X10Y7_E2BEG[7:0]),
	.E2BEGb(Tile_X10Y7_E2BEGb[7:0]),
	.EE4BEG(Tile_X10Y7_EE4BEG[15:0]),
	.E6BEG(Tile_X10Y7_E6BEG[11:0]),
	.S1BEG(Tile_X10Y7_S1BEG[3:0]),
	.S2BEG(Tile_X10Y7_S2BEG[7:0]),
	.S2BEGb(Tile_X10Y7_S2BEGb[7:0]),
	.S4BEG(Tile_X10Y7_S4BEG[15:0]),
	.SS4BEG(Tile_X10Y7_SS4BEG[15:0]),
	.W1BEG(Tile_X10Y7_W1BEG[3:0]),
	.W2BEG(Tile_X10Y7_W2BEG[7:0]),
	.W2BEGb(Tile_X10Y7_W2BEGb[7:0]),
	.WW4BEG(Tile_X10Y7_WW4BEG[15:0]),
	.W6BEG(Tile_X10Y7_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X10Y8_UserCLKo),
	.UserCLKo(Tile_X10Y7_UserCLKo),
	.FrameData(Tile_X9Y7_FrameData_O), 
	.FrameData_O(Tile_X10Y7_FrameData_O), 
	.FrameStrobe(Tile_X10Y8_FrameStrobe_O),
	.FrameStrobe_O(Tile_X10Y7_FrameStrobe_O)
	);

	E_CPU_IO Tile_X11Y7_E_CPU_IO (
	.E1END(Tile_X10Y7_E1BEG[3:0]),
	.E2MID(Tile_X10Y7_E2BEG[7:0]),
	.E2END(Tile_X10Y7_E2BEGb[7:0]),
	.EE4END(Tile_X10Y7_EE4BEG[15:0]),
	.E6END(Tile_X10Y7_E6BEG[11:0]),
	.W1BEG(Tile_X11Y7_W1BEG[3:0]),
	.W2BEG(Tile_X11Y7_W2BEG[7:0]),
	.W2BEGb(Tile_X11Y7_W2BEGb[7:0]),
	.WW4BEG(Tile_X11Y7_WW4BEG[15:0]),
	.W6BEG(Tile_X11Y7_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X11Y7_OPA_I0),
	.OPA_I1(Tile_X11Y7_OPA_I1),
	.OPA_I2(Tile_X11Y7_OPA_I2),
	.OPA_I3(Tile_X11Y7_OPA_I3),
	.UserCLK(Tile_X11Y8_UserCLKo),
	.OPB_I0(Tile_X11Y7_OPB_I0),
	.OPB_I1(Tile_X11Y7_OPB_I1),
	.OPB_I2(Tile_X11Y7_OPB_I2),
	.OPB_I3(Tile_X11Y7_OPB_I3),
	.RES0_O0(Tile_X11Y7_RES0_O0),
	.RES0_O1(Tile_X11Y7_RES0_O1),
	.RES0_O2(Tile_X11Y7_RES0_O2),
	.RES0_O3(Tile_X11Y7_RES0_O3),
	.RES1_O0(Tile_X11Y7_RES1_O0),
	.RES1_O1(Tile_X11Y7_RES1_O1),
	.RES1_O2(Tile_X11Y7_RES1_O2),
	.RES1_O3(Tile_X11Y7_RES1_O3),
	.RES2_O0(Tile_X11Y7_RES2_O0),
	.RES2_O1(Tile_X11Y7_RES2_O1),
	.RES2_O2(Tile_X11Y7_RES2_O2),
	.RES2_O3(Tile_X11Y7_RES2_O3),
	.UserCLKo(Tile_X11Y7_UserCLKo),
	.FrameData(Tile_X10Y7_FrameData_O), 
	.FrameData_O(Tile_X11Y7_FrameData_O), 
	.FrameStrobe(Tile_X11Y8_FrameStrobe_O),
	.FrameStrobe_O(Tile_X11Y7_FrameStrobe_O)
	);

	W_CPU_IO Tile_X4Y8_W_CPU_IO (
	.W1END(Tile_X5Y8_W1BEG[3:0]),
	.W2MID(Tile_X5Y8_W2BEG[7:0]),
	.W2END(Tile_X5Y8_W2BEGb[7:0]),
	.WW4END(Tile_X5Y8_WW4BEG[15:0]),
	.W6END(Tile_X5Y8_W6BEG[11:0]),
	.E1BEG(Tile_X4Y8_E1BEG[3:0]),
	.E2BEG(Tile_X4Y8_E2BEG[7:0]),
	.E2BEGb(Tile_X4Y8_E2BEGb[7:0]),
	.EE4BEG(Tile_X4Y8_EE4BEG[15:0]),
	.E6BEG(Tile_X4Y8_E6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X4Y8_OPA_I0),
	.OPA_I1(Tile_X4Y8_OPA_I1),
	.OPA_I2(Tile_X4Y8_OPA_I2),
	.OPA_I3(Tile_X4Y8_OPA_I3),
	.UserCLK(Tile_X4Y9_UserCLKo),
	.OPB_I0(Tile_X4Y8_OPB_I0),
	.OPB_I1(Tile_X4Y8_OPB_I1),
	.OPB_I2(Tile_X4Y8_OPB_I2),
	.OPB_I3(Tile_X4Y8_OPB_I3),
	.RES0_O0(Tile_X4Y8_RES0_O0),
	.RES0_O1(Tile_X4Y8_RES0_O1),
	.RES0_O2(Tile_X4Y8_RES0_O2),
	.RES0_O3(Tile_X4Y8_RES0_O3),
	.RES1_O0(Tile_X4Y8_RES1_O0),
	.RES1_O1(Tile_X4Y8_RES1_O1),
	.RES1_O2(Tile_X4Y8_RES1_O2),
	.RES1_O3(Tile_X4Y8_RES1_O3),
	.RES2_O0(Tile_X4Y8_RES2_O0),
	.RES2_O1(Tile_X4Y8_RES2_O1),
	.RES2_O2(Tile_X4Y8_RES2_O2),
	.RES2_O3(Tile_X4Y8_RES2_O3),
	.UserCLKo(Tile_X4Y8_UserCLKo),
	.FrameData(Tile_Y8_FrameData), 
	.FrameData_O(Tile_X4Y8_FrameData_O), 
	.FrameStrobe(Tile_X4Y9_FrameStrobe_O),
	.FrameStrobe_O(Tile_X4Y8_FrameStrobe_O)
	);


	LUT4AB Tile_X6Y8_LUT4AB (
	.N1END(Tile_X6Y9_N1BEG[3:0]),
	.N2MID(Tile_X6Y9_N2BEG[7:0]),
	.N2END(Tile_X6Y9_N2BEGb[7:0]),
	.N4END(Tile_X6Y9_N4BEG[15:0]),
	.NN4END(Tile_X6Y9_NN4BEG[15:0]),
	.Ci(Tile_X6Y9_Co[0:0]),
	.E1END(Tile_X5Y8_E1BEG[3:0]),
	.E2MID(Tile_X5Y8_E2BEG[7:0]),
	.E2END(Tile_X5Y8_E2BEGb[7:0]),
	.EE4END(Tile_X5Y8_EE4BEG[15:0]),
	.E6END(Tile_X5Y8_E6BEG[11:0]),
	.S1END(Tile_X6Y7_S1BEG[3:0]),
	.S2MID(Tile_X6Y7_S2BEG[7:0]),
	.S2END(Tile_X6Y7_S2BEGb[7:0]),
	.S4END(Tile_X6Y7_S4BEG[15:0]),
	.SS4END(Tile_X6Y7_SS4BEG[15:0]),
	.W1END(Tile_X7Y8_W1BEG[3:0]),
	.W2MID(Tile_X7Y8_W2BEG[7:0]),
	.W2END(Tile_X7Y8_W2BEGb[7:0]),
	.WW4END(Tile_X7Y8_WW4BEG[15:0]),
	.W6END(Tile_X7Y8_W6BEG[11:0]),
	.N1BEG(Tile_X6Y8_N1BEG[3:0]),
	.N2BEG(Tile_X6Y8_N2BEG[7:0]),
	.N2BEGb(Tile_X6Y8_N2BEGb[7:0]),
	.N4BEG(Tile_X6Y8_N4BEG[15:0]),
	.NN4BEG(Tile_X6Y8_NN4BEG[15:0]),
	.Co(Tile_X6Y8_Co[0:0]),
	.E1BEG(Tile_X6Y8_E1BEG[3:0]),
	.E2BEG(Tile_X6Y8_E2BEG[7:0]),
	.E2BEGb(Tile_X6Y8_E2BEGb[7:0]),
	.EE4BEG(Tile_X6Y8_EE4BEG[15:0]),
	.E6BEG(Tile_X6Y8_E6BEG[11:0]),
	.S1BEG(Tile_X6Y8_S1BEG[3:0]),
	.S2BEG(Tile_X6Y8_S2BEG[7:0]),
	.S2BEGb(Tile_X6Y8_S2BEGb[7:0]),
	.S4BEG(Tile_X6Y8_S4BEG[15:0]),
	.SS4BEG(Tile_X6Y8_SS4BEG[15:0]),
	.W1BEG(Tile_X6Y8_W1BEG[3:0]),
	.W2BEG(Tile_X6Y8_W2BEG[7:0]),
	.W2BEGb(Tile_X6Y8_W2BEGb[7:0]),
	.WW4BEG(Tile_X6Y8_WW4BEG[15:0]),
	.W6BEG(Tile_X6Y8_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X6Y9_UserCLKo),
	.UserCLKo(Tile_X6Y8_UserCLKo),
	.FrameData(Tile_X5Y8_FrameData_O), 
	.FrameData_O(Tile_X6Y8_FrameData_O), 
	.FrameStrobe(Tile_X6Y9_FrameStrobe_O),
	.FrameStrobe_O(Tile_X6Y8_FrameStrobe_O)
	);

	LUT4AB Tile_X7Y8_LUT4AB (
	.N1END(Tile_X7Y9_N1BEG[3:0]),
	.N2MID(Tile_X7Y9_N2BEG[7:0]),
	.N2END(Tile_X7Y9_N2BEGb[7:0]),
	.N4END(Tile_X7Y9_N4BEG[15:0]),
	.NN4END(Tile_X7Y9_NN4BEG[15:0]),
	.Ci(Tile_X7Y9_Co[0:0]),
	.E1END(Tile_X6Y8_E1BEG[3:0]),
	.E2MID(Tile_X6Y8_E2BEG[7:0]),
	.E2END(Tile_X6Y8_E2BEGb[7:0]),
	.EE4END(Tile_X6Y8_EE4BEG[15:0]),
	.E6END(Tile_X6Y8_E6BEG[11:0]),
	.S1END(Tile_X7Y7_S1BEG[3:0]),
	.S2MID(Tile_X7Y7_S2BEG[7:0]),
	.S2END(Tile_X7Y7_S2BEGb[7:0]),
	.S4END(Tile_X7Y7_S4BEG[15:0]),
	.SS4END(Tile_X7Y7_SS4BEG[15:0]),
	.W1END(Tile_X8Y8_W1BEG[3:0]),
	.W2MID(Tile_X8Y8_W2BEG[7:0]),
	.W2END(Tile_X8Y8_W2BEGb[7:0]),
	.WW4END(Tile_X8Y8_WW4BEG[15:0]),
	.W6END(Tile_X8Y8_W6BEG[11:0]),
	.N1BEG(Tile_X7Y8_N1BEG[3:0]),
	.N2BEG(Tile_X7Y8_N2BEG[7:0]),
	.N2BEGb(Tile_X7Y8_N2BEGb[7:0]),
	.N4BEG(Tile_X7Y8_N4BEG[15:0]),
	.NN4BEG(Tile_X7Y8_NN4BEG[15:0]),
	.Co(Tile_X7Y8_Co[0:0]),
	.E1BEG(Tile_X7Y8_E1BEG[3:0]),
	.E2BEG(Tile_X7Y8_E2BEG[7:0]),
	.E2BEGb(Tile_X7Y8_E2BEGb[7:0]),
	.EE4BEG(Tile_X7Y8_EE4BEG[15:0]),
	.E6BEG(Tile_X7Y8_E6BEG[11:0]),
	.S1BEG(Tile_X7Y8_S1BEG[3:0]),
	.S2BEG(Tile_X7Y8_S2BEG[7:0]),
	.S2BEGb(Tile_X7Y8_S2BEGb[7:0]),
	.S4BEG(Tile_X7Y8_S4BEG[15:0]),
	.SS4BEG(Tile_X7Y8_SS4BEG[15:0]),
	.W1BEG(Tile_X7Y8_W1BEG[3:0]),
	.W2BEG(Tile_X7Y8_W2BEG[7:0]),
	.W2BEGb(Tile_X7Y8_W2BEGb[7:0]),
	.WW4BEG(Tile_X7Y8_WW4BEG[15:0]),
	.W6BEG(Tile_X7Y8_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X7Y9_UserCLKo),
	.UserCLKo(Tile_X7Y8_UserCLKo),
	.FrameData(Tile_X6Y8_FrameData_O), 
	.FrameData_O(Tile_X7Y8_FrameData_O), 
	.FrameStrobe(Tile_X7Y9_FrameStrobe_O),
	.FrameStrobe_O(Tile_X7Y8_FrameStrobe_O)
	);

	LUT4AB Tile_X8Y8_LUT4AB (
	.N1END(Tile_X8Y9_N1BEG[3:0]),
	.N2MID(Tile_X8Y9_N2BEG[7:0]),
	.N2END(Tile_X8Y9_N2BEGb[7:0]),
	.N4END(Tile_X8Y9_N4BEG[15:0]),
	.NN4END(Tile_X8Y9_NN4BEG[15:0]),
	.Ci(Tile_X8Y9_Co[0:0]),
	.E1END(Tile_X7Y8_E1BEG[3:0]),
	.E2MID(Tile_X7Y8_E2BEG[7:0]),
	.E2END(Tile_X7Y8_E2BEGb[7:0]),
	.EE4END(Tile_X7Y8_EE4BEG[15:0]),
	.E6END(Tile_X7Y8_E6BEG[11:0]),
	.S1END(Tile_X8Y7_S1BEG[3:0]),
	.S2MID(Tile_X8Y7_S2BEG[7:0]),
	.S2END(Tile_X8Y7_S2BEGb[7:0]),
	.S4END(Tile_X8Y7_S4BEG[15:0]),
	.SS4END(Tile_X8Y7_SS4BEG[15:0]),
	.W1END(Tile_X9Y8_W1BEG[3:0]),
	.W2MID(Tile_X9Y8_W2BEG[7:0]),
	.W2END(Tile_X9Y8_W2BEGb[7:0]),
	.WW4END(Tile_X9Y8_WW4BEG[15:0]),
	.W6END(Tile_X9Y8_W6BEG[11:0]),
	.N1BEG(Tile_X8Y8_N1BEG[3:0]),
	.N2BEG(Tile_X8Y8_N2BEG[7:0]),
	.N2BEGb(Tile_X8Y8_N2BEGb[7:0]),
	.N4BEG(Tile_X8Y8_N4BEG[15:0]),
	.NN4BEG(Tile_X8Y8_NN4BEG[15:0]),
	.Co(Tile_X8Y8_Co[0:0]),
	.E1BEG(Tile_X8Y8_E1BEG[3:0]),
	.E2BEG(Tile_X8Y8_E2BEG[7:0]),
	.E2BEGb(Tile_X8Y8_E2BEGb[7:0]),
	.EE4BEG(Tile_X8Y8_EE4BEG[15:0]),
	.E6BEG(Tile_X8Y8_E6BEG[11:0]),
	.S1BEG(Tile_X8Y8_S1BEG[3:0]),
	.S2BEG(Tile_X8Y8_S2BEG[7:0]),
	.S2BEGb(Tile_X8Y8_S2BEGb[7:0]),
	.S4BEG(Tile_X8Y8_S4BEG[15:0]),
	.SS4BEG(Tile_X8Y8_SS4BEG[15:0]),
	.W1BEG(Tile_X8Y8_W1BEG[3:0]),
	.W2BEG(Tile_X8Y8_W2BEG[7:0]),
	.W2BEGb(Tile_X8Y8_W2BEGb[7:0]),
	.WW4BEG(Tile_X8Y8_WW4BEG[15:0]),
	.W6BEG(Tile_X8Y8_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X8Y9_UserCLKo),
	.UserCLKo(Tile_X8Y8_UserCLKo),
	.FrameData(Tile_X7Y8_FrameData_O), 
	.FrameData_O(Tile_X8Y8_FrameData_O), 
	.FrameStrobe(Tile_X8Y9_FrameStrobe_O),
	.FrameStrobe_O(Tile_X8Y8_FrameStrobe_O)
	);


	LUT4AB Tile_X10Y8_LUT4AB (
	.N1END(Tile_X10Y9_N1BEG[3:0]),
	.N2MID(Tile_X10Y9_N2BEG[7:0]),
	.N2END(Tile_X10Y9_N2BEGb[7:0]),
	.N4END(Tile_X10Y9_N4BEG[15:0]),
	.NN4END(Tile_X10Y9_NN4BEG[15:0]),
	.Ci(Tile_X10Y9_Co[0:0]),
	.E1END(Tile_X9Y8_E1BEG[3:0]),
	.E2MID(Tile_X9Y8_E2BEG[7:0]),
	.E2END(Tile_X9Y8_E2BEGb[7:0]),
	.EE4END(Tile_X9Y8_EE4BEG[15:0]),
	.E6END(Tile_X9Y8_E6BEG[11:0]),
	.S1END(Tile_X10Y7_S1BEG[3:0]),
	.S2MID(Tile_X10Y7_S2BEG[7:0]),
	.S2END(Tile_X10Y7_S2BEGb[7:0]),
	.S4END(Tile_X10Y7_S4BEG[15:0]),
	.SS4END(Tile_X10Y7_SS4BEG[15:0]),
	.W1END(Tile_X11Y8_W1BEG[3:0]),
	.W2MID(Tile_X11Y8_W2BEG[7:0]),
	.W2END(Tile_X11Y8_W2BEGb[7:0]),
	.WW4END(Tile_X11Y8_WW4BEG[15:0]),
	.W6END(Tile_X11Y8_W6BEG[11:0]),
	.N1BEG(Tile_X10Y8_N1BEG[3:0]),
	.N2BEG(Tile_X10Y8_N2BEG[7:0]),
	.N2BEGb(Tile_X10Y8_N2BEGb[7:0]),
	.N4BEG(Tile_X10Y8_N4BEG[15:0]),
	.NN4BEG(Tile_X10Y8_NN4BEG[15:0]),
	.Co(Tile_X10Y8_Co[0:0]),
	.E1BEG(Tile_X10Y8_E1BEG[3:0]),
	.E2BEG(Tile_X10Y8_E2BEG[7:0]),
	.E2BEGb(Tile_X10Y8_E2BEGb[7:0]),
	.EE4BEG(Tile_X10Y8_EE4BEG[15:0]),
	.E6BEG(Tile_X10Y8_E6BEG[11:0]),
	.S1BEG(Tile_X10Y8_S1BEG[3:0]),
	.S2BEG(Tile_X10Y8_S2BEG[7:0]),
	.S2BEGb(Tile_X10Y8_S2BEGb[7:0]),
	.S4BEG(Tile_X10Y8_S4BEG[15:0]),
	.SS4BEG(Tile_X10Y8_SS4BEG[15:0]),
	.W1BEG(Tile_X10Y8_W1BEG[3:0]),
	.W2BEG(Tile_X10Y8_W2BEG[7:0]),
	.W2BEGb(Tile_X10Y8_W2BEGb[7:0]),
	.WW4BEG(Tile_X10Y8_WW4BEG[15:0]),
	.W6BEG(Tile_X10Y8_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X10Y9_UserCLKo),
	.UserCLKo(Tile_X10Y8_UserCLKo),
	.FrameData(Tile_X9Y8_FrameData_O), 
	.FrameData_O(Tile_X10Y8_FrameData_O), 
	.FrameStrobe(Tile_X10Y9_FrameStrobe_O),
	.FrameStrobe_O(Tile_X10Y8_FrameStrobe_O)
	);

	E_CPU_IO Tile_X11Y8_E_CPU_IO (
	.E1END(Tile_X10Y8_E1BEG[3:0]),
	.E2MID(Tile_X10Y8_E2BEG[7:0]),
	.E2END(Tile_X10Y8_E2BEGb[7:0]),
	.EE4END(Tile_X10Y8_EE4BEG[15:0]),
	.E6END(Tile_X10Y8_E6BEG[11:0]),
	.W1BEG(Tile_X11Y8_W1BEG[3:0]),
	.W2BEG(Tile_X11Y8_W2BEG[7:0]),
	.W2BEGb(Tile_X11Y8_W2BEGb[7:0]),
	.WW4BEG(Tile_X11Y8_WW4BEG[15:0]),
	.W6BEG(Tile_X11Y8_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X11Y8_OPA_I0),
	.OPA_I1(Tile_X11Y8_OPA_I1),
	.OPA_I2(Tile_X11Y8_OPA_I2),
	.OPA_I3(Tile_X11Y8_OPA_I3),
	.UserCLK(Tile_X11Y9_UserCLKo),
	.OPB_I0(Tile_X11Y8_OPB_I0),
	.OPB_I1(Tile_X11Y8_OPB_I1),
	.OPB_I2(Tile_X11Y8_OPB_I2),
	.OPB_I3(Tile_X11Y8_OPB_I3),
	.RES0_O0(Tile_X11Y8_RES0_O0),
	.RES0_O1(Tile_X11Y8_RES0_O1),
	.RES0_O2(Tile_X11Y8_RES0_O2),
	.RES0_O3(Tile_X11Y8_RES0_O3),
	.RES1_O0(Tile_X11Y8_RES1_O0),
	.RES1_O1(Tile_X11Y8_RES1_O1),
	.RES1_O2(Tile_X11Y8_RES1_O2),
	.RES1_O3(Tile_X11Y8_RES1_O3),
	.RES2_O0(Tile_X11Y8_RES2_O0),
	.RES2_O1(Tile_X11Y8_RES2_O1),
	.RES2_O2(Tile_X11Y8_RES2_O2),
	.RES2_O3(Tile_X11Y8_RES2_O3),
	.UserCLKo(Tile_X11Y8_UserCLKo),
	.FrameData(Tile_X10Y8_FrameData_O), 
	.FrameData_O(Tile_X11Y8_FrameData_O), 
	.FrameStrobe(Tile_X11Y9_FrameStrobe_O),
	.FrameStrobe_O(Tile_X11Y8_FrameStrobe_O)
	);

	N_term_single Tile_X1Y9_N_term_single (
	.N1END(Tile_X1Y10_N1BEG[3:0]),
	.N2MID(Tile_X1Y10_N2BEG[7:0]),
	.N2END(Tile_X1Y10_N2BEGb[7:0]),
	.N4END(Tile_X1Y10_N4BEG[15:0]),
	.NN4END(Tile_X1Y10_NN4BEG[15:0]),
	.Ci(Tile_X1Y10_Co[0:0]),
	.S1BEG(Tile_X1Y9_S1BEG[3:0]),
	.S2BEG(Tile_X1Y9_S2BEG[7:0]),
	.S2BEGb(Tile_X1Y9_S2BEGb[7:0]),
	.S4BEG(Tile_X1Y9_S4BEG[15:0]),
	.SS4BEG(Tile_X1Y9_SS4BEG[15:0]),
	.UserCLK(Tile_X1Y10_UserCLKo),
	.UserCLKo(Tile_X1Y9_UserCLKo),
	.FrameStrobe(Tile_X1Y10_FrameStrobe_O),
	.FrameStrobe_O(Tile_X1Y9_FrameStrobe_O)
	);

	N_term_single2 Tile_X2Y9_N_term_single2 (
	.N1END(Tile_X2Y10_N1BEG[3:0]),
	.N2MID(Tile_X2Y10_N2BEG[7:0]),
	.N2END(Tile_X2Y10_N2BEGb[7:0]),
	.N4END(Tile_X2Y10_N4BEG[15:0]),
	.NN4END(Tile_X2Y10_NN4BEG[15:0]),
	.S1BEG(Tile_X2Y9_S1BEG[3:0]),
	.S2BEG(Tile_X2Y9_S2BEG[7:0]),
	.S2BEGb(Tile_X2Y9_S2BEGb[7:0]),
	.S4BEG(Tile_X2Y9_S4BEG[15:0]),
	.SS4BEG(Tile_X2Y9_SS4BEG[15:0]),
	.UserCLK(Tile_X2Y10_UserCLKo),
	.UserCLKo(Tile_X2Y9_UserCLKo),
	.FrameStrobe(Tile_X2Y10_FrameStrobe_O),
	.FrameStrobe_O(Tile_X2Y9_FrameStrobe_O)
	);

	N_term_single Tile_X3Y9_N_term_single (
	.N1END(Tile_X3Y10_N1BEG[3:0]),
	.N2MID(Tile_X3Y10_N2BEG[7:0]),
	.N2END(Tile_X3Y10_N2BEGb[7:0]),
	.N4END(Tile_X3Y10_N4BEG[15:0]),
	.NN4END(Tile_X3Y10_NN4BEG[15:0]),
	.Ci(Tile_X3Y10_Co[0:0]),
	.S1BEG(Tile_X3Y9_S1BEG[3:0]),
	.S2BEG(Tile_X3Y9_S2BEG[7:0]),
	.S2BEGb(Tile_X3Y9_S2BEGb[7:0]),
	.S4BEG(Tile_X3Y9_S4BEG[15:0]),
	.SS4BEG(Tile_X3Y9_SS4BEG[15:0]),
	.UserCLK(Tile_X3Y10_UserCLKo),
	.UserCLKo(Tile_X3Y9_UserCLKo),
	.FrameStrobe(Tile_X3Y10_FrameStrobe_O),
	.FrameStrobe_O(Tile_X3Y9_FrameStrobe_O)
	);

	W_CPU_IO_bot Tile_X4Y9_W_CPU_IO_bot (
	.N1END(Tile_X4Y10_N1BEG[3:0]),
	.N2MID(Tile_X4Y10_N2BEG[7:0]),
	.N2END(Tile_X4Y10_N2BEGb[7:0]),
	.N4END(Tile_X4Y10_N4BEG[15:0]),
	.NN4END(Tile_X4Y10_NN4BEG[15:0]),
	.Ci(Tile_X4Y10_Co[0:0]),
	.W1END(Tile_X5Y9_W1BEG[3:0]),
	.W2MID(Tile_X5Y9_W2BEG[7:0]),
	.W2END(Tile_X5Y9_W2BEGb[7:0]),
	.WW4END(Tile_X5Y9_WW4BEG[15:0]),
	.W6END(Tile_X5Y9_W6BEG[11:0]),
	.E1BEG(Tile_X4Y9_E1BEG[3:0]),
	.E2BEG(Tile_X4Y9_E2BEG[7:0]),
	.E2BEGb(Tile_X4Y9_E2BEGb[7:0]),
	.EE4BEG(Tile_X4Y9_EE4BEG[15:0]),
	.E6BEG(Tile_X4Y9_E6BEG[11:0]),
	.S1BEG(Tile_X4Y9_S1BEG[3:0]),
	.S2BEG(Tile_X4Y9_S2BEG[7:0]),
	.S2BEGb(Tile_X4Y9_S2BEGb[7:0]),
	.S4BEG(Tile_X4Y9_S4BEG[15:0]),
	.SS4BEG(Tile_X4Y9_SS4BEG[15:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X4Y9_OPA_I0),
	.OPA_I1(Tile_X4Y9_OPA_I1),
	.OPA_I2(Tile_X4Y9_OPA_I2),
	.OPA_I3(Tile_X4Y9_OPA_I3),
	.UserCLK(Tile_X4Y10_UserCLKo),
	.OPB_I0(Tile_X4Y9_OPB_I0),
	.OPB_I1(Tile_X4Y9_OPB_I1),
	.OPB_I2(Tile_X4Y9_OPB_I2),
	.OPB_I3(Tile_X4Y9_OPB_I3),
	.RES0_O0(Tile_X4Y9_RES0_O0),
	.RES0_O1(Tile_X4Y9_RES0_O1),
	.RES0_O2(Tile_X4Y9_RES0_O2),
	.RES0_O3(Tile_X4Y9_RES0_O3),
	.RES1_O0(Tile_X4Y9_RES1_O0),
	.RES1_O1(Tile_X4Y9_RES1_O1),
	.RES1_O2(Tile_X4Y9_RES1_O2),
	.RES1_O3(Tile_X4Y9_RES1_O3),
	.RES2_O0(Tile_X4Y9_RES2_O0),
	.RES2_O1(Tile_X4Y9_RES2_O1),
	.RES2_O2(Tile_X4Y9_RES2_O2),
	.RES2_O3(Tile_X4Y9_RES2_O3),
	.UserCLKo(Tile_X4Y9_UserCLKo),
	.FrameData(Tile_Y9_FrameData), 
	.FrameData_O(Tile_X4Y9_FrameData_O), 
	.FrameStrobe(Tile_X4Y10_FrameStrobe_O),
	.FrameStrobe_O(Tile_X4Y9_FrameStrobe_O)
	);


	LUT4AB Tile_X6Y9_LUT4AB (
	.N1END(Tile_X6Y10_N1BEG[3:0]),
	.N2MID(Tile_X6Y10_N2BEG[7:0]),
	.N2END(Tile_X6Y10_N2BEGb[7:0]),
	.N4END(Tile_X6Y10_N4BEG[15:0]),
	.NN4END(Tile_X6Y10_NN4BEG[15:0]),
	.Ci(Tile_X6Y10_Co[0:0]),
	.E1END(Tile_X5Y9_E1BEG[3:0]),
	.E2MID(Tile_X5Y9_E2BEG[7:0]),
	.E2END(Tile_X5Y9_E2BEGb[7:0]),
	.EE4END(Tile_X5Y9_EE4BEG[15:0]),
	.E6END(Tile_X5Y9_E6BEG[11:0]),
	.S1END(Tile_X6Y8_S1BEG[3:0]),
	.S2MID(Tile_X6Y8_S2BEG[7:0]),
	.S2END(Tile_X6Y8_S2BEGb[7:0]),
	.S4END(Tile_X6Y8_S4BEG[15:0]),
	.SS4END(Tile_X6Y8_SS4BEG[15:0]),
	.W1END(Tile_X7Y9_W1BEG[3:0]),
	.W2MID(Tile_X7Y9_W2BEG[7:0]),
	.W2END(Tile_X7Y9_W2BEGb[7:0]),
	.WW4END(Tile_X7Y9_WW4BEG[15:0]),
	.W6END(Tile_X7Y9_W6BEG[11:0]),
	.N1BEG(Tile_X6Y9_N1BEG[3:0]),
	.N2BEG(Tile_X6Y9_N2BEG[7:0]),
	.N2BEGb(Tile_X6Y9_N2BEGb[7:0]),
	.N4BEG(Tile_X6Y9_N4BEG[15:0]),
	.NN4BEG(Tile_X6Y9_NN4BEG[15:0]),
	.Co(Tile_X6Y9_Co[0:0]),
	.E1BEG(Tile_X6Y9_E1BEG[3:0]),
	.E2BEG(Tile_X6Y9_E2BEG[7:0]),
	.E2BEGb(Tile_X6Y9_E2BEGb[7:0]),
	.EE4BEG(Tile_X6Y9_EE4BEG[15:0]),
	.E6BEG(Tile_X6Y9_E6BEG[11:0]),
	.S1BEG(Tile_X6Y9_S1BEG[3:0]),
	.S2BEG(Tile_X6Y9_S2BEG[7:0]),
	.S2BEGb(Tile_X6Y9_S2BEGb[7:0]),
	.S4BEG(Tile_X6Y9_S4BEG[15:0]),
	.SS4BEG(Tile_X6Y9_SS4BEG[15:0]),
	.W1BEG(Tile_X6Y9_W1BEG[3:0]),
	.W2BEG(Tile_X6Y9_W2BEG[7:0]),
	.W2BEGb(Tile_X6Y9_W2BEGb[7:0]),
	.WW4BEG(Tile_X6Y9_WW4BEG[15:0]),
	.W6BEG(Tile_X6Y9_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X6Y10_UserCLKo),
	.UserCLKo(Tile_X6Y9_UserCLKo),
	.FrameData(Tile_X5Y9_FrameData_O), 
	.FrameData_O(Tile_X6Y9_FrameData_O), 
	.FrameStrobe(Tile_X6Y10_FrameStrobe_O),
	.FrameStrobe_O(Tile_X6Y9_FrameStrobe_O)
	);

	LUT4AB Tile_X7Y9_LUT4AB (
	.N1END(Tile_X7Y10_N1BEG[3:0]),
	.N2MID(Tile_X7Y10_N2BEG[7:0]),
	.N2END(Tile_X7Y10_N2BEGb[7:0]),
	.N4END(Tile_X7Y10_N4BEG[15:0]),
	.NN4END(Tile_X7Y10_NN4BEG[15:0]),
	.Ci(Tile_X7Y10_Co[0:0]),
	.E1END(Tile_X6Y9_E1BEG[3:0]),
	.E2MID(Tile_X6Y9_E2BEG[7:0]),
	.E2END(Tile_X6Y9_E2BEGb[7:0]),
	.EE4END(Tile_X6Y9_EE4BEG[15:0]),
	.E6END(Tile_X6Y9_E6BEG[11:0]),
	.S1END(Tile_X7Y8_S1BEG[3:0]),
	.S2MID(Tile_X7Y8_S2BEG[7:0]),
	.S2END(Tile_X7Y8_S2BEGb[7:0]),
	.S4END(Tile_X7Y8_S4BEG[15:0]),
	.SS4END(Tile_X7Y8_SS4BEG[15:0]),
	.W1END(Tile_X8Y9_W1BEG[3:0]),
	.W2MID(Tile_X8Y9_W2BEG[7:0]),
	.W2END(Tile_X8Y9_W2BEGb[7:0]),
	.WW4END(Tile_X8Y9_WW4BEG[15:0]),
	.W6END(Tile_X8Y9_W6BEG[11:0]),
	.N1BEG(Tile_X7Y9_N1BEG[3:0]),
	.N2BEG(Tile_X7Y9_N2BEG[7:0]),
	.N2BEGb(Tile_X7Y9_N2BEGb[7:0]),
	.N4BEG(Tile_X7Y9_N4BEG[15:0]),
	.NN4BEG(Tile_X7Y9_NN4BEG[15:0]),
	.Co(Tile_X7Y9_Co[0:0]),
	.E1BEG(Tile_X7Y9_E1BEG[3:0]),
	.E2BEG(Tile_X7Y9_E2BEG[7:0]),
	.E2BEGb(Tile_X7Y9_E2BEGb[7:0]),
	.EE4BEG(Tile_X7Y9_EE4BEG[15:0]),
	.E6BEG(Tile_X7Y9_E6BEG[11:0]),
	.S1BEG(Tile_X7Y9_S1BEG[3:0]),
	.S2BEG(Tile_X7Y9_S2BEG[7:0]),
	.S2BEGb(Tile_X7Y9_S2BEGb[7:0]),
	.S4BEG(Tile_X7Y9_S4BEG[15:0]),
	.SS4BEG(Tile_X7Y9_SS4BEG[15:0]),
	.W1BEG(Tile_X7Y9_W1BEG[3:0]),
	.W2BEG(Tile_X7Y9_W2BEG[7:0]),
	.W2BEGb(Tile_X7Y9_W2BEGb[7:0]),
	.WW4BEG(Tile_X7Y9_WW4BEG[15:0]),
	.W6BEG(Tile_X7Y9_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X7Y10_UserCLKo),
	.UserCLKo(Tile_X7Y9_UserCLKo),
	.FrameData(Tile_X6Y9_FrameData_O), 
	.FrameData_O(Tile_X7Y9_FrameData_O), 
	.FrameStrobe(Tile_X7Y10_FrameStrobe_O),
	.FrameStrobe_O(Tile_X7Y9_FrameStrobe_O)
	);

	LUT4AB Tile_X8Y9_LUT4AB (
	.N1END(Tile_X8Y10_N1BEG[3:0]),
	.N2MID(Tile_X8Y10_N2BEG[7:0]),
	.N2END(Tile_X8Y10_N2BEGb[7:0]),
	.N4END(Tile_X8Y10_N4BEG[15:0]),
	.NN4END(Tile_X8Y10_NN4BEG[15:0]),
	.Ci(Tile_X8Y10_Co[0:0]),
	.E1END(Tile_X7Y9_E1BEG[3:0]),
	.E2MID(Tile_X7Y9_E2BEG[7:0]),
	.E2END(Tile_X7Y9_E2BEGb[7:0]),
	.EE4END(Tile_X7Y9_EE4BEG[15:0]),
	.E6END(Tile_X7Y9_E6BEG[11:0]),
	.S1END(Tile_X8Y8_S1BEG[3:0]),
	.S2MID(Tile_X8Y8_S2BEG[7:0]),
	.S2END(Tile_X8Y8_S2BEGb[7:0]),
	.S4END(Tile_X8Y8_S4BEG[15:0]),
	.SS4END(Tile_X8Y8_SS4BEG[15:0]),
	.W1END(Tile_X9Y9_W1BEG[3:0]),
	.W2MID(Tile_X9Y9_W2BEG[7:0]),
	.W2END(Tile_X9Y9_W2BEGb[7:0]),
	.WW4END(Tile_X9Y9_WW4BEG[15:0]),
	.W6END(Tile_X9Y9_W6BEG[11:0]),
	.N1BEG(Tile_X8Y9_N1BEG[3:0]),
	.N2BEG(Tile_X8Y9_N2BEG[7:0]),
	.N2BEGb(Tile_X8Y9_N2BEGb[7:0]),
	.N4BEG(Tile_X8Y9_N4BEG[15:0]),
	.NN4BEG(Tile_X8Y9_NN4BEG[15:0]),
	.Co(Tile_X8Y9_Co[0:0]),
	.E1BEG(Tile_X8Y9_E1BEG[3:0]),
	.E2BEG(Tile_X8Y9_E2BEG[7:0]),
	.E2BEGb(Tile_X8Y9_E2BEGb[7:0]),
	.EE4BEG(Tile_X8Y9_EE4BEG[15:0]),
	.E6BEG(Tile_X8Y9_E6BEG[11:0]),
	.S1BEG(Tile_X8Y9_S1BEG[3:0]),
	.S2BEG(Tile_X8Y9_S2BEG[7:0]),
	.S2BEGb(Tile_X8Y9_S2BEGb[7:0]),
	.S4BEG(Tile_X8Y9_S4BEG[15:0]),
	.SS4BEG(Tile_X8Y9_SS4BEG[15:0]),
	.W1BEG(Tile_X8Y9_W1BEG[3:0]),
	.W2BEG(Tile_X8Y9_W2BEG[7:0]),
	.W2BEGb(Tile_X8Y9_W2BEGb[7:0]),
	.WW4BEG(Tile_X8Y9_WW4BEG[15:0]),
	.W6BEG(Tile_X8Y9_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X8Y10_UserCLKo),
	.UserCLKo(Tile_X8Y9_UserCLKo),
	.FrameData(Tile_X7Y9_FrameData_O), 
	.FrameData_O(Tile_X8Y9_FrameData_O), 
	.FrameStrobe(Tile_X8Y10_FrameStrobe_O),
	.FrameStrobe_O(Tile_X8Y9_FrameStrobe_O)
	);


	LUT4AB Tile_X10Y9_LUT4AB (
	.N1END(Tile_X10Y10_N1BEG[3:0]),
	.N2MID(Tile_X10Y10_N2BEG[7:0]),
	.N2END(Tile_X10Y10_N2BEGb[7:0]),
	.N4END(Tile_X10Y10_N4BEG[15:0]),
	.NN4END(Tile_X10Y10_NN4BEG[15:0]),
	.Ci(Tile_X10Y10_Co[0:0]),
	.E1END(Tile_X9Y9_E1BEG[3:0]),
	.E2MID(Tile_X9Y9_E2BEG[7:0]),
	.E2END(Tile_X9Y9_E2BEGb[7:0]),
	.EE4END(Tile_X9Y9_EE4BEG[15:0]),
	.E6END(Tile_X9Y9_E6BEG[11:0]),
	.S1END(Tile_X10Y8_S1BEG[3:0]),
	.S2MID(Tile_X10Y8_S2BEG[7:0]),
	.S2END(Tile_X10Y8_S2BEGb[7:0]),
	.S4END(Tile_X10Y8_S4BEG[15:0]),
	.SS4END(Tile_X10Y8_SS4BEG[15:0]),
	.W1END(Tile_X11Y9_W1BEG[3:0]),
	.W2MID(Tile_X11Y9_W2BEG[7:0]),
	.W2END(Tile_X11Y9_W2BEGb[7:0]),
	.WW4END(Tile_X11Y9_WW4BEG[15:0]),
	.W6END(Tile_X11Y9_W6BEG[11:0]),
	.N1BEG(Tile_X10Y9_N1BEG[3:0]),
	.N2BEG(Tile_X10Y9_N2BEG[7:0]),
	.N2BEGb(Tile_X10Y9_N2BEGb[7:0]),
	.N4BEG(Tile_X10Y9_N4BEG[15:0]),
	.NN4BEG(Tile_X10Y9_NN4BEG[15:0]),
	.Co(Tile_X10Y9_Co[0:0]),
	.E1BEG(Tile_X10Y9_E1BEG[3:0]),
	.E2BEG(Tile_X10Y9_E2BEG[7:0]),
	.E2BEGb(Tile_X10Y9_E2BEGb[7:0]),
	.EE4BEG(Tile_X10Y9_EE4BEG[15:0]),
	.E6BEG(Tile_X10Y9_E6BEG[11:0]),
	.S1BEG(Tile_X10Y9_S1BEG[3:0]),
	.S2BEG(Tile_X10Y9_S2BEG[7:0]),
	.S2BEGb(Tile_X10Y9_S2BEGb[7:0]),
	.S4BEG(Tile_X10Y9_S4BEG[15:0]),
	.SS4BEG(Tile_X10Y9_SS4BEG[15:0]),
	.W1BEG(Tile_X10Y9_W1BEG[3:0]),
	.W2BEG(Tile_X10Y9_W2BEG[7:0]),
	.W2BEGb(Tile_X10Y9_W2BEGb[7:0]),
	.WW4BEG(Tile_X10Y9_WW4BEG[15:0]),
	.W6BEG(Tile_X10Y9_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X10Y10_UserCLKo),
	.UserCLKo(Tile_X10Y9_UserCLKo),
	.FrameData(Tile_X9Y9_FrameData_O), 
	.FrameData_O(Tile_X10Y9_FrameData_O), 
	.FrameStrobe(Tile_X10Y10_FrameStrobe_O),
	.FrameStrobe_O(Tile_X10Y9_FrameStrobe_O)
	);

	E_CPU_IO_bot Tile_X11Y9_E_CPU_IO_bot (
	.N1END(Tile_X11Y10_N1BEG[3:0]),
	.N2MID(Tile_X11Y10_N2BEG[7:0]),
	.N2END(Tile_X11Y10_N2BEGb[7:0]),
	.N4END(Tile_X11Y10_N4BEG[15:0]),
	.NN4END(Tile_X11Y10_NN4BEG[15:0]),
	.Ci(Tile_X11Y10_Co[0:0]),
	.E1END(Tile_X10Y9_E1BEG[3:0]),
	.E2MID(Tile_X10Y9_E2BEG[7:0]),
	.E2END(Tile_X10Y9_E2BEGb[7:0]),
	.EE4END(Tile_X10Y9_EE4BEG[15:0]),
	.E6END(Tile_X10Y9_E6BEG[11:0]),
	.S1BEG(Tile_X11Y9_S1BEG[3:0]),
	.S2BEG(Tile_X11Y9_S2BEG[7:0]),
	.S2BEGb(Tile_X11Y9_S2BEGb[7:0]),
	.S4BEG(Tile_X11Y9_S4BEG[15:0]),
	.SS4BEG(Tile_X11Y9_SS4BEG[15:0]),
	.W1BEG(Tile_X11Y9_W1BEG[3:0]),
	.W2BEG(Tile_X11Y9_W2BEG[7:0]),
	.W2BEGb(Tile_X11Y9_W2BEGb[7:0]),
	.WW4BEG(Tile_X11Y9_WW4BEG[15:0]),
	.W6BEG(Tile_X11Y9_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X11Y9_OPA_I0),
	.OPA_I1(Tile_X11Y9_OPA_I1),
	.OPA_I2(Tile_X11Y9_OPA_I2),
	.OPA_I3(Tile_X11Y9_OPA_I3),
	.UserCLK(Tile_X11Y10_UserCLKo),
	.OPB_I0(Tile_X11Y9_OPB_I0),
	.OPB_I1(Tile_X11Y9_OPB_I1),
	.OPB_I2(Tile_X11Y9_OPB_I2),
	.OPB_I3(Tile_X11Y9_OPB_I3),
	.RES0_O0(Tile_X11Y9_RES0_O0),
	.RES0_O1(Tile_X11Y9_RES0_O1),
	.RES0_O2(Tile_X11Y9_RES0_O2),
	.RES0_O3(Tile_X11Y9_RES0_O3),
	.RES1_O0(Tile_X11Y9_RES1_O0),
	.RES1_O1(Tile_X11Y9_RES1_O1),
	.RES1_O2(Tile_X11Y9_RES1_O2),
	.RES1_O3(Tile_X11Y9_RES1_O3),
	.RES2_O0(Tile_X11Y9_RES2_O0),
	.RES2_O1(Tile_X11Y9_RES2_O1),
	.RES2_O2(Tile_X11Y9_RES2_O2),
	.RES2_O3(Tile_X11Y9_RES2_O3),
	.UserCLKo(Tile_X11Y9_UserCLKo),
	.FrameData(Tile_X10Y9_FrameData_O), 
	.FrameData_O(Tile_X11Y9_FrameData_O), 
	.FrameStrobe(Tile_X11Y10_FrameStrobe_O),
	.FrameStrobe_O(Tile_X11Y9_FrameStrobe_O)
	);

	N_term_single Tile_X12Y9_N_term_single (
	.N1END(Tile_X12Y10_N1BEG[3:0]),
	.N2MID(Tile_X12Y10_N2BEG[7:0]),
	.N2END(Tile_X12Y10_N2BEGb[7:0]),
	.N4END(Tile_X12Y10_N4BEG[15:0]),
	.NN4END(Tile_X12Y10_NN4BEG[15:0]),
	.Ci(Tile_X12Y10_Co[0:0]),
	.S1BEG(Tile_X12Y9_S1BEG[3:0]),
	.S2BEG(Tile_X12Y9_S2BEG[7:0]),
	.S2BEGb(Tile_X12Y9_S2BEGb[7:0]),
	.S4BEG(Tile_X12Y9_S4BEG[15:0]),
	.SS4BEG(Tile_X12Y9_SS4BEG[15:0]),
	.UserCLK(Tile_X12Y10_UserCLKo),
	.UserCLKo(Tile_X12Y9_UserCLKo),
	.FrameStrobe(Tile_X12Y10_FrameStrobe_O),
	.FrameStrobe_O(Tile_X12Y9_FrameStrobe_O)
	);

	N_term_single2 Tile_X13Y9_N_term_single2 (
	.N1END(Tile_X13Y10_N1BEG[3:0]),
	.N2MID(Tile_X13Y10_N2BEG[7:0]),
	.N2END(Tile_X13Y10_N2BEGb[7:0]),
	.N4END(Tile_X13Y10_N4BEG[15:0]),
	.NN4END(Tile_X13Y10_NN4BEG[15:0]),
	.S1BEG(Tile_X13Y9_S1BEG[3:0]),
	.S2BEG(Tile_X13Y9_S2BEG[7:0]),
	.S2BEGb(Tile_X13Y9_S2BEGb[7:0]),
	.S4BEG(Tile_X13Y9_S4BEG[15:0]),
	.SS4BEG(Tile_X13Y9_SS4BEG[15:0]),
	.UserCLK(Tile_X13Y10_UserCLKo),
	.UserCLKo(Tile_X13Y9_UserCLKo),
	.FrameStrobe(Tile_X13Y10_FrameStrobe_O),
	.FrameStrobe_O(Tile_X13Y9_FrameStrobe_O)
	);

	N_term_single Tile_X14Y9_N_term_single (
	.N1END(Tile_X14Y10_N1BEG[3:0]),
	.N2MID(Tile_X14Y10_N2BEG[7:0]),
	.N2END(Tile_X14Y10_N2BEGb[7:0]),
	.N4END(Tile_X14Y10_N4BEG[15:0]),
	.NN4END(Tile_X14Y10_NN4BEG[15:0]),
	.Ci(Tile_X14Y10_Co[0:0]),
	.S1BEG(Tile_X14Y9_S1BEG[3:0]),
	.S2BEG(Tile_X14Y9_S2BEG[7:0]),
	.S2BEGb(Tile_X14Y9_S2BEGb[7:0]),
	.S4BEG(Tile_X14Y9_S4BEG[15:0]),
	.SS4BEG(Tile_X14Y9_SS4BEG[15:0]),
	.UserCLK(Tile_X14Y10_UserCLKo),
	.UserCLKo(Tile_X14Y9_UserCLKo),
	.FrameStrobe(Tile_X14Y10_FrameStrobe_O),
	.FrameStrobe_O(Tile_X14Y9_FrameStrobe_O)
	);

	N_term_RAM_IO Tile_X15Y9_N_term_RAM_IO (
	.N1END(Tile_X15Y10_N1BEG[3:0]),
	.N2MID(Tile_X15Y10_N2BEG[7:0]),
	.N2END(Tile_X15Y10_N2BEGb[7:0]),
	.N4END(Tile_X15Y10_N4BEG[15:0]),
	.S1BEG(Tile_X15Y9_S1BEG[3:0]),
	.S2BEG(Tile_X15Y9_S2BEG[7:0]),
	.S2BEGb(Tile_X15Y9_S2BEGb[7:0]),
	.S4BEG(Tile_X15Y9_S4BEG[15:0]),
	.UserCLK(Tile_X15Y10_UserCLKo),
	.UserCLKo(Tile_X15Y9_UserCLKo),
	.FrameStrobe(Tile_X15Y10_FrameStrobe_O),
	.FrameStrobe_O(Tile_X15Y9_FrameStrobe_O)
	);

	W_IO Tile_X0Y10_W_IO (
	.W1END(Tile_X1Y10_W1BEG[3:0]),
	.W2MID(Tile_X1Y10_W2BEG[7:0]),
	.W2END(Tile_X1Y10_W2BEGb[7:0]),
	.WW4END(Tile_X1Y10_WW4BEG[15:0]),
	.W6END(Tile_X1Y10_W6BEG[11:0]),
	.E1BEG(Tile_X0Y10_E1BEG[3:0]),
	.E2BEG(Tile_X0Y10_E2BEG[7:0]),
	.E2BEGb(Tile_X0Y10_E2BEGb[7:0]),
	.EE4BEG(Tile_X0Y10_EE4BEG[15:0]),
	.E6BEG(Tile_X0Y10_E6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.A_I_top(Tile_X0Y10_A_I_top),
	.A_T_top(Tile_X0Y10_A_T_top),
	.A_O_top(Tile_X0Y10_A_O_top),
	.UserCLK(Tile_X0Y11_UserCLKo),
	.B_I_top(Tile_X0Y10_B_I_top),
	.B_T_top(Tile_X0Y10_B_T_top),
	.B_O_top(Tile_X0Y10_B_O_top),
	.A_config_C_bit0(Tile_X0Y10_A_config_C_bit0),
	.A_config_C_bit1(Tile_X0Y10_A_config_C_bit1),
	.A_config_C_bit2(Tile_X0Y10_A_config_C_bit2),
	.A_config_C_bit3(Tile_X0Y10_A_config_C_bit3),
	.B_config_C_bit0(Tile_X0Y10_B_config_C_bit0),
	.B_config_C_bit1(Tile_X0Y10_B_config_C_bit1),
	.B_config_C_bit2(Tile_X0Y10_B_config_C_bit2),
	.B_config_C_bit3(Tile_X0Y10_B_config_C_bit3),
	.UserCLKo(Tile_X0Y10_UserCLKo),
	.FrameData(Tile_Y10_FrameData), 
	.FrameData_O(Tile_X0Y10_FrameData_O), 
	.FrameStrobe(Tile_X0Y11_FrameStrobe_O),
	.FrameStrobe_O(Tile_X0Y10_FrameStrobe_O)
	);

	LUT4AB Tile_X1Y10_LUT4AB (
	.N1END(Tile_X1Y11_N1BEG[3:0]),
	.N2MID(Tile_X1Y11_N2BEG[7:0]),
	.N2END(Tile_X1Y11_N2BEGb[7:0]),
	.N4END(Tile_X1Y11_N4BEG[15:0]),
	.NN4END(Tile_X1Y11_NN4BEG[15:0]),
	.Ci(Tile_X1Y11_Co[0:0]),
	.E1END(Tile_X0Y10_E1BEG[3:0]),
	.E2MID(Tile_X0Y10_E2BEG[7:0]),
	.E2END(Tile_X0Y10_E2BEGb[7:0]),
	.EE4END(Tile_X0Y10_EE4BEG[15:0]),
	.E6END(Tile_X0Y10_E6BEG[11:0]),
	.S1END(Tile_X1Y9_S1BEG[3:0]),
	.S2MID(Tile_X1Y9_S2BEG[7:0]),
	.S2END(Tile_X1Y9_S2BEGb[7:0]),
	.S4END(Tile_X1Y9_S4BEG[15:0]),
	.SS4END(Tile_X1Y9_SS4BEG[15:0]),
	.W1END(Tile_X2Y10_W1BEG[3:0]),
	.W2MID(Tile_X2Y10_W2BEG[7:0]),
	.W2END(Tile_X2Y10_W2BEGb[7:0]),
	.WW4END(Tile_X2Y10_WW4BEG[15:0]),
	.W6END(Tile_X2Y10_W6BEG[11:0]),
	.N1BEG(Tile_X1Y10_N1BEG[3:0]),
	.N2BEG(Tile_X1Y10_N2BEG[7:0]),
	.N2BEGb(Tile_X1Y10_N2BEGb[7:0]),
	.N4BEG(Tile_X1Y10_N4BEG[15:0]),
	.NN4BEG(Tile_X1Y10_NN4BEG[15:0]),
	.Co(Tile_X1Y10_Co[0:0]),
	.E1BEG(Tile_X1Y10_E1BEG[3:0]),
	.E2BEG(Tile_X1Y10_E2BEG[7:0]),
	.E2BEGb(Tile_X1Y10_E2BEGb[7:0]),
	.EE4BEG(Tile_X1Y10_EE4BEG[15:0]),
	.E6BEG(Tile_X1Y10_E6BEG[11:0]),
	.S1BEG(Tile_X1Y10_S1BEG[3:0]),
	.S2BEG(Tile_X1Y10_S2BEG[7:0]),
	.S2BEGb(Tile_X1Y10_S2BEGb[7:0]),
	.S4BEG(Tile_X1Y10_S4BEG[15:0]),
	.SS4BEG(Tile_X1Y10_SS4BEG[15:0]),
	.W1BEG(Tile_X1Y10_W1BEG[3:0]),
	.W2BEG(Tile_X1Y10_W2BEG[7:0]),
	.W2BEGb(Tile_X1Y10_W2BEGb[7:0]),
	.WW4BEG(Tile_X1Y10_WW4BEG[15:0]),
	.W6BEG(Tile_X1Y10_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X1Y11_UserCLKo),
	.UserCLKo(Tile_X1Y10_UserCLKo),
	.FrameData(Tile_X0Y10_FrameData_O), 
	.FrameData_O(Tile_X1Y10_FrameData_O), 
	.FrameStrobe(Tile_X1Y11_FrameStrobe_O),
	.FrameStrobe_O(Tile_X1Y10_FrameStrobe_O)
	);

	RegFile Tile_X2Y10_RegFile (
	.N1END(Tile_X2Y11_N1BEG[3:0]),
	.N2MID(Tile_X2Y11_N2BEG[7:0]),
	.N2END(Tile_X2Y11_N2BEGb[7:0]),
	.N4END(Tile_X2Y11_N4BEG[15:0]),
	.NN4END(Tile_X2Y11_NN4BEG[15:0]),
	.E1END(Tile_X1Y10_E1BEG[3:0]),
	.E2MID(Tile_X1Y10_E2BEG[7:0]),
	.E2END(Tile_X1Y10_E2BEGb[7:0]),
	.EE4END(Tile_X1Y10_EE4BEG[15:0]),
	.E6END(Tile_X1Y10_E6BEG[11:0]),
	.S1END(Tile_X2Y9_S1BEG[3:0]),
	.S2MID(Tile_X2Y9_S2BEG[7:0]),
	.S2END(Tile_X2Y9_S2BEGb[7:0]),
	.S4END(Tile_X2Y9_S4BEG[15:0]),
	.SS4END(Tile_X2Y9_SS4BEG[15:0]),
	.W1END(Tile_X3Y10_W1BEG[3:0]),
	.W2MID(Tile_X3Y10_W2BEG[7:0]),
	.W2END(Tile_X3Y10_W2BEGb[7:0]),
	.WW4END(Tile_X3Y10_WW4BEG[15:0]),
	.W6END(Tile_X3Y10_W6BEG[11:0]),
	.N1BEG(Tile_X2Y10_N1BEG[3:0]),
	.N2BEG(Tile_X2Y10_N2BEG[7:0]),
	.N2BEGb(Tile_X2Y10_N2BEGb[7:0]),
	.N4BEG(Tile_X2Y10_N4BEG[15:0]),
	.NN4BEG(Tile_X2Y10_NN4BEG[15:0]),
	.E1BEG(Tile_X2Y10_E1BEG[3:0]),
	.E2BEG(Tile_X2Y10_E2BEG[7:0]),
	.E2BEGb(Tile_X2Y10_E2BEGb[7:0]),
	.EE4BEG(Tile_X2Y10_EE4BEG[15:0]),
	.E6BEG(Tile_X2Y10_E6BEG[11:0]),
	.S1BEG(Tile_X2Y10_S1BEG[3:0]),
	.S2BEG(Tile_X2Y10_S2BEG[7:0]),
	.S2BEGb(Tile_X2Y10_S2BEGb[7:0]),
	.S4BEG(Tile_X2Y10_S4BEG[15:0]),
	.SS4BEG(Tile_X2Y10_SS4BEG[15:0]),
	.W1BEG(Tile_X2Y10_W1BEG[3:0]),
	.W2BEG(Tile_X2Y10_W2BEG[7:0]),
	.W2BEGb(Tile_X2Y10_W2BEGb[7:0]),
	.WW4BEG(Tile_X2Y10_WW4BEG[15:0]),
	.W6BEG(Tile_X2Y10_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X2Y11_UserCLKo),
	.UserCLKo(Tile_X2Y10_UserCLKo),
	.FrameData(Tile_X1Y10_FrameData_O), 
	.FrameData_O(Tile_X2Y10_FrameData_O), 
	.FrameStrobe(Tile_X2Y11_FrameStrobe_O),
	.FrameStrobe_O(Tile_X2Y10_FrameStrobe_O)
	);

	LUT4AB Tile_X3Y10_LUT4AB (
	.N1END(Tile_X3Y11_N1BEG[3:0]),
	.N2MID(Tile_X3Y11_N2BEG[7:0]),
	.N2END(Tile_X3Y11_N2BEGb[7:0]),
	.N4END(Tile_X3Y11_N4BEG[15:0]),
	.NN4END(Tile_X3Y11_NN4BEG[15:0]),
	.Ci(Tile_X3Y11_Co[0:0]),
	.E1END(Tile_X2Y10_E1BEG[3:0]),
	.E2MID(Tile_X2Y10_E2BEG[7:0]),
	.E2END(Tile_X2Y10_E2BEGb[7:0]),
	.EE4END(Tile_X2Y10_EE4BEG[15:0]),
	.E6END(Tile_X2Y10_E6BEG[11:0]),
	.S1END(Tile_X3Y9_S1BEG[3:0]),
	.S2MID(Tile_X3Y9_S2BEG[7:0]),
	.S2END(Tile_X3Y9_S2BEGb[7:0]),
	.S4END(Tile_X3Y9_S4BEG[15:0]),
	.SS4END(Tile_X3Y9_SS4BEG[15:0]),
	.W1END(Tile_X4Y10_W1BEG[3:0]),
	.W2MID(Tile_X4Y10_W2BEG[7:0]),
	.W2END(Tile_X4Y10_W2BEGb[7:0]),
	.WW4END(Tile_X4Y10_WW4BEG[15:0]),
	.W6END(Tile_X4Y10_W6BEG[11:0]),
	.N1BEG(Tile_X3Y10_N1BEG[3:0]),
	.N2BEG(Tile_X3Y10_N2BEG[7:0]),
	.N2BEGb(Tile_X3Y10_N2BEGb[7:0]),
	.N4BEG(Tile_X3Y10_N4BEG[15:0]),
	.NN4BEG(Tile_X3Y10_NN4BEG[15:0]),
	.Co(Tile_X3Y10_Co[0:0]),
	.E1BEG(Tile_X3Y10_E1BEG[3:0]),
	.E2BEG(Tile_X3Y10_E2BEG[7:0]),
	.E2BEGb(Tile_X3Y10_E2BEGb[7:0]),
	.EE4BEG(Tile_X3Y10_EE4BEG[15:0]),
	.E6BEG(Tile_X3Y10_E6BEG[11:0]),
	.S1BEG(Tile_X3Y10_S1BEG[3:0]),
	.S2BEG(Tile_X3Y10_S2BEG[7:0]),
	.S2BEGb(Tile_X3Y10_S2BEGb[7:0]),
	.S4BEG(Tile_X3Y10_S4BEG[15:0]),
	.SS4BEG(Tile_X3Y10_SS4BEG[15:0]),
	.W1BEG(Tile_X3Y10_W1BEG[3:0]),
	.W2BEG(Tile_X3Y10_W2BEG[7:0]),
	.W2BEGb(Tile_X3Y10_W2BEGb[7:0]),
	.WW4BEG(Tile_X3Y10_WW4BEG[15:0]),
	.W6BEG(Tile_X3Y10_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X3Y11_UserCLKo),
	.UserCLKo(Tile_X3Y10_UserCLKo),
	.FrameData(Tile_X2Y10_FrameData_O), 
	.FrameData_O(Tile_X3Y10_FrameData_O), 
	.FrameStrobe(Tile_X3Y11_FrameStrobe_O),
	.FrameStrobe_O(Tile_X3Y10_FrameStrobe_O)
	);

	LUT4AB Tile_X4Y10_LUT4AB (
	.N1END(Tile_X4Y11_N1BEG[3:0]),
	.N2MID(Tile_X4Y11_N2BEG[7:0]),
	.N2END(Tile_X4Y11_N2BEGb[7:0]),
	.N4END(Tile_X4Y11_N4BEG[15:0]),
	.NN4END(Tile_X4Y11_NN4BEG[15:0]),
	.Ci(Tile_X4Y11_Co[0:0]),
	.E1END(Tile_X3Y10_E1BEG[3:0]),
	.E2MID(Tile_X3Y10_E2BEG[7:0]),
	.E2END(Tile_X3Y10_E2BEGb[7:0]),
	.EE4END(Tile_X3Y10_EE4BEG[15:0]),
	.E6END(Tile_X3Y10_E6BEG[11:0]),
	.S1END(Tile_X4Y9_S1BEG[3:0]),
	.S2MID(Tile_X4Y9_S2BEG[7:0]),
	.S2END(Tile_X4Y9_S2BEGb[7:0]),
	.S4END(Tile_X4Y9_S4BEG[15:0]),
	.SS4END(Tile_X4Y9_SS4BEG[15:0]),
	.W1END(Tile_X5Y10_W1BEG[3:0]),
	.W2MID(Tile_X5Y10_W2BEG[7:0]),
	.W2END(Tile_X5Y10_W2BEGb[7:0]),
	.WW4END(Tile_X5Y10_WW4BEG[15:0]),
	.W6END(Tile_X5Y10_W6BEG[11:0]),
	.N1BEG(Tile_X4Y10_N1BEG[3:0]),
	.N2BEG(Tile_X4Y10_N2BEG[7:0]),
	.N2BEGb(Tile_X4Y10_N2BEGb[7:0]),
	.N4BEG(Tile_X4Y10_N4BEG[15:0]),
	.NN4BEG(Tile_X4Y10_NN4BEG[15:0]),
	.Co(Tile_X4Y10_Co[0:0]),
	.E1BEG(Tile_X4Y10_E1BEG[3:0]),
	.E2BEG(Tile_X4Y10_E2BEG[7:0]),
	.E2BEGb(Tile_X4Y10_E2BEGb[7:0]),
	.EE4BEG(Tile_X4Y10_EE4BEG[15:0]),
	.E6BEG(Tile_X4Y10_E6BEG[11:0]),
	.S1BEG(Tile_X4Y10_S1BEG[3:0]),
	.S2BEG(Tile_X4Y10_S2BEG[7:0]),
	.S2BEGb(Tile_X4Y10_S2BEGb[7:0]),
	.S4BEG(Tile_X4Y10_S4BEG[15:0]),
	.SS4BEG(Tile_X4Y10_SS4BEG[15:0]),
	.W1BEG(Tile_X4Y10_W1BEG[3:0]),
	.W2BEG(Tile_X4Y10_W2BEG[7:0]),
	.W2BEGb(Tile_X4Y10_W2BEGb[7:0]),
	.WW4BEG(Tile_X4Y10_WW4BEG[15:0]),
	.W6BEG(Tile_X4Y10_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X4Y11_UserCLKo),
	.UserCLKo(Tile_X4Y10_UserCLKo),
	.FrameData(Tile_X3Y10_FrameData_O), 
	.FrameData_O(Tile_X4Y10_FrameData_O), 
	.FrameStrobe(Tile_X4Y11_FrameStrobe_O),
	.FrameStrobe_O(Tile_X4Y10_FrameStrobe_O)
	);


	LUT4AB Tile_X6Y10_LUT4AB (
	.N1END(Tile_X6Y11_N1BEG[3:0]),
	.N2MID(Tile_X6Y11_N2BEG[7:0]),
	.N2END(Tile_X6Y11_N2BEGb[7:0]),
	.N4END(Tile_X6Y11_N4BEG[15:0]),
	.NN4END(Tile_X6Y11_NN4BEG[15:0]),
	.Ci(Tile_X6Y11_Co[0:0]),
	.E1END(Tile_X5Y10_E1BEG[3:0]),
	.E2MID(Tile_X5Y10_E2BEG[7:0]),
	.E2END(Tile_X5Y10_E2BEGb[7:0]),
	.EE4END(Tile_X5Y10_EE4BEG[15:0]),
	.E6END(Tile_X5Y10_E6BEG[11:0]),
	.S1END(Tile_X6Y9_S1BEG[3:0]),
	.S2MID(Tile_X6Y9_S2BEG[7:0]),
	.S2END(Tile_X6Y9_S2BEGb[7:0]),
	.S4END(Tile_X6Y9_S4BEG[15:0]),
	.SS4END(Tile_X6Y9_SS4BEG[15:0]),
	.W1END(Tile_X7Y10_W1BEG[3:0]),
	.W2MID(Tile_X7Y10_W2BEG[7:0]),
	.W2END(Tile_X7Y10_W2BEGb[7:0]),
	.WW4END(Tile_X7Y10_WW4BEG[15:0]),
	.W6END(Tile_X7Y10_W6BEG[11:0]),
	.N1BEG(Tile_X6Y10_N1BEG[3:0]),
	.N2BEG(Tile_X6Y10_N2BEG[7:0]),
	.N2BEGb(Tile_X6Y10_N2BEGb[7:0]),
	.N4BEG(Tile_X6Y10_N4BEG[15:0]),
	.NN4BEG(Tile_X6Y10_NN4BEG[15:0]),
	.Co(Tile_X6Y10_Co[0:0]),
	.E1BEG(Tile_X6Y10_E1BEG[3:0]),
	.E2BEG(Tile_X6Y10_E2BEG[7:0]),
	.E2BEGb(Tile_X6Y10_E2BEGb[7:0]),
	.EE4BEG(Tile_X6Y10_EE4BEG[15:0]),
	.E6BEG(Tile_X6Y10_E6BEG[11:0]),
	.S1BEG(Tile_X6Y10_S1BEG[3:0]),
	.S2BEG(Tile_X6Y10_S2BEG[7:0]),
	.S2BEGb(Tile_X6Y10_S2BEGb[7:0]),
	.S4BEG(Tile_X6Y10_S4BEG[15:0]),
	.SS4BEG(Tile_X6Y10_SS4BEG[15:0]),
	.W1BEG(Tile_X6Y10_W1BEG[3:0]),
	.W2BEG(Tile_X6Y10_W2BEG[7:0]),
	.W2BEGb(Tile_X6Y10_W2BEGb[7:0]),
	.WW4BEG(Tile_X6Y10_WW4BEG[15:0]),
	.W6BEG(Tile_X6Y10_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X6Y11_UserCLKo),
	.UserCLKo(Tile_X6Y10_UserCLKo),
	.FrameData(Tile_X5Y10_FrameData_O), 
	.FrameData_O(Tile_X6Y10_FrameData_O), 
	.FrameStrobe(Tile_X6Y11_FrameStrobe_O),
	.FrameStrobe_O(Tile_X6Y10_FrameStrobe_O)
	);

	LUT4AB Tile_X7Y10_LUT4AB (
	.N1END(Tile_X7Y11_N1BEG[3:0]),
	.N2MID(Tile_X7Y11_N2BEG[7:0]),
	.N2END(Tile_X7Y11_N2BEGb[7:0]),
	.N4END(Tile_X7Y11_N4BEG[15:0]),
	.NN4END(Tile_X7Y11_NN4BEG[15:0]),
	.Ci(Tile_X7Y11_Co[0:0]),
	.E1END(Tile_X6Y10_E1BEG[3:0]),
	.E2MID(Tile_X6Y10_E2BEG[7:0]),
	.E2END(Tile_X6Y10_E2BEGb[7:0]),
	.EE4END(Tile_X6Y10_EE4BEG[15:0]),
	.E6END(Tile_X6Y10_E6BEG[11:0]),
	.S1END(Tile_X7Y9_S1BEG[3:0]),
	.S2MID(Tile_X7Y9_S2BEG[7:0]),
	.S2END(Tile_X7Y9_S2BEGb[7:0]),
	.S4END(Tile_X7Y9_S4BEG[15:0]),
	.SS4END(Tile_X7Y9_SS4BEG[15:0]),
	.W1END(Tile_X8Y10_W1BEG[3:0]),
	.W2MID(Tile_X8Y10_W2BEG[7:0]),
	.W2END(Tile_X8Y10_W2BEGb[7:0]),
	.WW4END(Tile_X8Y10_WW4BEG[15:0]),
	.W6END(Tile_X8Y10_W6BEG[11:0]),
	.N1BEG(Tile_X7Y10_N1BEG[3:0]),
	.N2BEG(Tile_X7Y10_N2BEG[7:0]),
	.N2BEGb(Tile_X7Y10_N2BEGb[7:0]),
	.N4BEG(Tile_X7Y10_N4BEG[15:0]),
	.NN4BEG(Tile_X7Y10_NN4BEG[15:0]),
	.Co(Tile_X7Y10_Co[0:0]),
	.E1BEG(Tile_X7Y10_E1BEG[3:0]),
	.E2BEG(Tile_X7Y10_E2BEG[7:0]),
	.E2BEGb(Tile_X7Y10_E2BEGb[7:0]),
	.EE4BEG(Tile_X7Y10_EE4BEG[15:0]),
	.E6BEG(Tile_X7Y10_E6BEG[11:0]),
	.S1BEG(Tile_X7Y10_S1BEG[3:0]),
	.S2BEG(Tile_X7Y10_S2BEG[7:0]),
	.S2BEGb(Tile_X7Y10_S2BEGb[7:0]),
	.S4BEG(Tile_X7Y10_S4BEG[15:0]),
	.SS4BEG(Tile_X7Y10_SS4BEG[15:0]),
	.W1BEG(Tile_X7Y10_W1BEG[3:0]),
	.W2BEG(Tile_X7Y10_W2BEG[7:0]),
	.W2BEGb(Tile_X7Y10_W2BEGb[7:0]),
	.WW4BEG(Tile_X7Y10_WW4BEG[15:0]),
	.W6BEG(Tile_X7Y10_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X7Y11_UserCLKo),
	.UserCLKo(Tile_X7Y10_UserCLKo),
	.FrameData(Tile_X6Y10_FrameData_O), 
	.FrameData_O(Tile_X7Y10_FrameData_O), 
	.FrameStrobe(Tile_X7Y11_FrameStrobe_O),
	.FrameStrobe_O(Tile_X7Y10_FrameStrobe_O)
	);

	LUT4AB Tile_X8Y10_LUT4AB (
	.N1END(Tile_X8Y11_N1BEG[3:0]),
	.N2MID(Tile_X8Y11_N2BEG[7:0]),
	.N2END(Tile_X8Y11_N2BEGb[7:0]),
	.N4END(Tile_X8Y11_N4BEG[15:0]),
	.NN4END(Tile_X8Y11_NN4BEG[15:0]),
	.Ci(Tile_X8Y11_Co[0:0]),
	.E1END(Tile_X7Y10_E1BEG[3:0]),
	.E2MID(Tile_X7Y10_E2BEG[7:0]),
	.E2END(Tile_X7Y10_E2BEGb[7:0]),
	.EE4END(Tile_X7Y10_EE4BEG[15:0]),
	.E6END(Tile_X7Y10_E6BEG[11:0]),
	.S1END(Tile_X8Y9_S1BEG[3:0]),
	.S2MID(Tile_X8Y9_S2BEG[7:0]),
	.S2END(Tile_X8Y9_S2BEGb[7:0]),
	.S4END(Tile_X8Y9_S4BEG[15:0]),
	.SS4END(Tile_X8Y9_SS4BEG[15:0]),
	.W1END(Tile_X9Y10_W1BEG[3:0]),
	.W2MID(Tile_X9Y10_W2BEG[7:0]),
	.W2END(Tile_X9Y10_W2BEGb[7:0]),
	.WW4END(Tile_X9Y10_WW4BEG[15:0]),
	.W6END(Tile_X9Y10_W6BEG[11:0]),
	.N1BEG(Tile_X8Y10_N1BEG[3:0]),
	.N2BEG(Tile_X8Y10_N2BEG[7:0]),
	.N2BEGb(Tile_X8Y10_N2BEGb[7:0]),
	.N4BEG(Tile_X8Y10_N4BEG[15:0]),
	.NN4BEG(Tile_X8Y10_NN4BEG[15:0]),
	.Co(Tile_X8Y10_Co[0:0]),
	.E1BEG(Tile_X8Y10_E1BEG[3:0]),
	.E2BEG(Tile_X8Y10_E2BEG[7:0]),
	.E2BEGb(Tile_X8Y10_E2BEGb[7:0]),
	.EE4BEG(Tile_X8Y10_EE4BEG[15:0]),
	.E6BEG(Tile_X8Y10_E6BEG[11:0]),
	.S1BEG(Tile_X8Y10_S1BEG[3:0]),
	.S2BEG(Tile_X8Y10_S2BEG[7:0]),
	.S2BEGb(Tile_X8Y10_S2BEGb[7:0]),
	.S4BEG(Tile_X8Y10_S4BEG[15:0]),
	.SS4BEG(Tile_X8Y10_SS4BEG[15:0]),
	.W1BEG(Tile_X8Y10_W1BEG[3:0]),
	.W2BEG(Tile_X8Y10_W2BEG[7:0]),
	.W2BEGb(Tile_X8Y10_W2BEGb[7:0]),
	.WW4BEG(Tile_X8Y10_WW4BEG[15:0]),
	.W6BEG(Tile_X8Y10_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X8Y11_UserCLKo),
	.UserCLKo(Tile_X8Y10_UserCLKo),
	.FrameData(Tile_X7Y10_FrameData_O), 
	.FrameData_O(Tile_X8Y10_FrameData_O), 
	.FrameStrobe(Tile_X8Y11_FrameStrobe_O),
	.FrameStrobe_O(Tile_X8Y10_FrameStrobe_O)
	);


	LUT4AB Tile_X10Y10_LUT4AB (
	.N1END(Tile_X10Y11_N1BEG[3:0]),
	.N2MID(Tile_X10Y11_N2BEG[7:0]),
	.N2END(Tile_X10Y11_N2BEGb[7:0]),
	.N4END(Tile_X10Y11_N4BEG[15:0]),
	.NN4END(Tile_X10Y11_NN4BEG[15:0]),
	.Ci(Tile_X10Y11_Co[0:0]),
	.E1END(Tile_X9Y10_E1BEG[3:0]),
	.E2MID(Tile_X9Y10_E2BEG[7:0]),
	.E2END(Tile_X9Y10_E2BEGb[7:0]),
	.EE4END(Tile_X9Y10_EE4BEG[15:0]),
	.E6END(Tile_X9Y10_E6BEG[11:0]),
	.S1END(Tile_X10Y9_S1BEG[3:0]),
	.S2MID(Tile_X10Y9_S2BEG[7:0]),
	.S2END(Tile_X10Y9_S2BEGb[7:0]),
	.S4END(Tile_X10Y9_S4BEG[15:0]),
	.SS4END(Tile_X10Y9_SS4BEG[15:0]),
	.W1END(Tile_X11Y10_W1BEG[3:0]),
	.W2MID(Tile_X11Y10_W2BEG[7:0]),
	.W2END(Tile_X11Y10_W2BEGb[7:0]),
	.WW4END(Tile_X11Y10_WW4BEG[15:0]),
	.W6END(Tile_X11Y10_W6BEG[11:0]),
	.N1BEG(Tile_X10Y10_N1BEG[3:0]),
	.N2BEG(Tile_X10Y10_N2BEG[7:0]),
	.N2BEGb(Tile_X10Y10_N2BEGb[7:0]),
	.N4BEG(Tile_X10Y10_N4BEG[15:0]),
	.NN4BEG(Tile_X10Y10_NN4BEG[15:0]),
	.Co(Tile_X10Y10_Co[0:0]),
	.E1BEG(Tile_X10Y10_E1BEG[3:0]),
	.E2BEG(Tile_X10Y10_E2BEG[7:0]),
	.E2BEGb(Tile_X10Y10_E2BEGb[7:0]),
	.EE4BEG(Tile_X10Y10_EE4BEG[15:0]),
	.E6BEG(Tile_X10Y10_E6BEG[11:0]),
	.S1BEG(Tile_X10Y10_S1BEG[3:0]),
	.S2BEG(Tile_X10Y10_S2BEG[7:0]),
	.S2BEGb(Tile_X10Y10_S2BEGb[7:0]),
	.S4BEG(Tile_X10Y10_S4BEG[15:0]),
	.SS4BEG(Tile_X10Y10_SS4BEG[15:0]),
	.W1BEG(Tile_X10Y10_W1BEG[3:0]),
	.W2BEG(Tile_X10Y10_W2BEG[7:0]),
	.W2BEGb(Tile_X10Y10_W2BEGb[7:0]),
	.WW4BEG(Tile_X10Y10_WW4BEG[15:0]),
	.W6BEG(Tile_X10Y10_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X10Y11_UserCLKo),
	.UserCLKo(Tile_X10Y10_UserCLKo),
	.FrameData(Tile_X9Y10_FrameData_O), 
	.FrameData_O(Tile_X10Y10_FrameData_O), 
	.FrameStrobe(Tile_X10Y11_FrameStrobe_O),
	.FrameStrobe_O(Tile_X10Y10_FrameStrobe_O)
	);

	LUT4AB Tile_X11Y10_LUT4AB (
	.N1END(Tile_X11Y11_N1BEG[3:0]),
	.N2MID(Tile_X11Y11_N2BEG[7:0]),
	.N2END(Tile_X11Y11_N2BEGb[7:0]),
	.N4END(Tile_X11Y11_N4BEG[15:0]),
	.NN4END(Tile_X11Y11_NN4BEG[15:0]),
	.Ci(Tile_X11Y11_Co[0:0]),
	.E1END(Tile_X10Y10_E1BEG[3:0]),
	.E2MID(Tile_X10Y10_E2BEG[7:0]),
	.E2END(Tile_X10Y10_E2BEGb[7:0]),
	.EE4END(Tile_X10Y10_EE4BEG[15:0]),
	.E6END(Tile_X10Y10_E6BEG[11:0]),
	.S1END(Tile_X11Y9_S1BEG[3:0]),
	.S2MID(Tile_X11Y9_S2BEG[7:0]),
	.S2END(Tile_X11Y9_S2BEGb[7:0]),
	.S4END(Tile_X11Y9_S4BEG[15:0]),
	.SS4END(Tile_X11Y9_SS4BEG[15:0]),
	.W1END(Tile_X12Y10_W1BEG[3:0]),
	.W2MID(Tile_X12Y10_W2BEG[7:0]),
	.W2END(Tile_X12Y10_W2BEGb[7:0]),
	.WW4END(Tile_X12Y10_WW4BEG[15:0]),
	.W6END(Tile_X12Y10_W6BEG[11:0]),
	.N1BEG(Tile_X11Y10_N1BEG[3:0]),
	.N2BEG(Tile_X11Y10_N2BEG[7:0]),
	.N2BEGb(Tile_X11Y10_N2BEGb[7:0]),
	.N4BEG(Tile_X11Y10_N4BEG[15:0]),
	.NN4BEG(Tile_X11Y10_NN4BEG[15:0]),
	.Co(Tile_X11Y10_Co[0:0]),
	.E1BEG(Tile_X11Y10_E1BEG[3:0]),
	.E2BEG(Tile_X11Y10_E2BEG[7:0]),
	.E2BEGb(Tile_X11Y10_E2BEGb[7:0]),
	.EE4BEG(Tile_X11Y10_EE4BEG[15:0]),
	.E6BEG(Tile_X11Y10_E6BEG[11:0]),
	.S1BEG(Tile_X11Y10_S1BEG[3:0]),
	.S2BEG(Tile_X11Y10_S2BEG[7:0]),
	.S2BEGb(Tile_X11Y10_S2BEGb[7:0]),
	.S4BEG(Tile_X11Y10_S4BEG[15:0]),
	.SS4BEG(Tile_X11Y10_SS4BEG[15:0]),
	.W1BEG(Tile_X11Y10_W1BEG[3:0]),
	.W2BEG(Tile_X11Y10_W2BEG[7:0]),
	.W2BEGb(Tile_X11Y10_W2BEGb[7:0]),
	.WW4BEG(Tile_X11Y10_WW4BEG[15:0]),
	.W6BEG(Tile_X11Y10_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X11Y11_UserCLKo),
	.UserCLKo(Tile_X11Y10_UserCLKo),
	.FrameData(Tile_X10Y10_FrameData_O), 
	.FrameData_O(Tile_X11Y10_FrameData_O), 
	.FrameStrobe(Tile_X11Y11_FrameStrobe_O),
	.FrameStrobe_O(Tile_X11Y10_FrameStrobe_O)
	);

	LUT4AB Tile_X12Y10_LUT4AB (
	.N1END(Tile_X12Y11_N1BEG[3:0]),
	.N2MID(Tile_X12Y11_N2BEG[7:0]),
	.N2END(Tile_X12Y11_N2BEGb[7:0]),
	.N4END(Tile_X12Y11_N4BEG[15:0]),
	.NN4END(Tile_X12Y11_NN4BEG[15:0]),
	.Ci(Tile_X12Y11_Co[0:0]),
	.E1END(Tile_X11Y10_E1BEG[3:0]),
	.E2MID(Tile_X11Y10_E2BEG[7:0]),
	.E2END(Tile_X11Y10_E2BEGb[7:0]),
	.EE4END(Tile_X11Y10_EE4BEG[15:0]),
	.E6END(Tile_X11Y10_E6BEG[11:0]),
	.S1END(Tile_X12Y9_S1BEG[3:0]),
	.S2MID(Tile_X12Y9_S2BEG[7:0]),
	.S2END(Tile_X12Y9_S2BEGb[7:0]),
	.S4END(Tile_X12Y9_S4BEG[15:0]),
	.SS4END(Tile_X12Y9_SS4BEG[15:0]),
	.W1END(Tile_X13Y10_W1BEG[3:0]),
	.W2MID(Tile_X13Y10_W2BEG[7:0]),
	.W2END(Tile_X13Y10_W2BEGb[7:0]),
	.WW4END(Tile_X13Y10_WW4BEG[15:0]),
	.W6END(Tile_X13Y10_W6BEG[11:0]),
	.N1BEG(Tile_X12Y10_N1BEG[3:0]),
	.N2BEG(Tile_X12Y10_N2BEG[7:0]),
	.N2BEGb(Tile_X12Y10_N2BEGb[7:0]),
	.N4BEG(Tile_X12Y10_N4BEG[15:0]),
	.NN4BEG(Tile_X12Y10_NN4BEG[15:0]),
	.Co(Tile_X12Y10_Co[0:0]),
	.E1BEG(Tile_X12Y10_E1BEG[3:0]),
	.E2BEG(Tile_X12Y10_E2BEG[7:0]),
	.E2BEGb(Tile_X12Y10_E2BEGb[7:0]),
	.EE4BEG(Tile_X12Y10_EE4BEG[15:0]),
	.E6BEG(Tile_X12Y10_E6BEG[11:0]),
	.S1BEG(Tile_X12Y10_S1BEG[3:0]),
	.S2BEG(Tile_X12Y10_S2BEG[7:0]),
	.S2BEGb(Tile_X12Y10_S2BEGb[7:0]),
	.S4BEG(Tile_X12Y10_S4BEG[15:0]),
	.SS4BEG(Tile_X12Y10_SS4BEG[15:0]),
	.W1BEG(Tile_X12Y10_W1BEG[3:0]),
	.W2BEG(Tile_X12Y10_W2BEG[7:0]),
	.W2BEGb(Tile_X12Y10_W2BEGb[7:0]),
	.WW4BEG(Tile_X12Y10_WW4BEG[15:0]),
	.W6BEG(Tile_X12Y10_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X12Y11_UserCLKo),
	.UserCLKo(Tile_X12Y10_UserCLKo),
	.FrameData(Tile_X11Y10_FrameData_O), 
	.FrameData_O(Tile_X12Y10_FrameData_O), 
	.FrameStrobe(Tile_X12Y11_FrameStrobe_O),
	.FrameStrobe_O(Tile_X12Y10_FrameStrobe_O)
	);

	RegFile Tile_X13Y10_RegFile (
	.N1END(Tile_X13Y11_N1BEG[3:0]),
	.N2MID(Tile_X13Y11_N2BEG[7:0]),
	.N2END(Tile_X13Y11_N2BEGb[7:0]),
	.N4END(Tile_X13Y11_N4BEG[15:0]),
	.NN4END(Tile_X13Y11_NN4BEG[15:0]),
	.E1END(Tile_X12Y10_E1BEG[3:0]),
	.E2MID(Tile_X12Y10_E2BEG[7:0]),
	.E2END(Tile_X12Y10_E2BEGb[7:0]),
	.EE4END(Tile_X12Y10_EE4BEG[15:0]),
	.E6END(Tile_X12Y10_E6BEG[11:0]),
	.S1END(Tile_X13Y9_S1BEG[3:0]),
	.S2MID(Tile_X13Y9_S2BEG[7:0]),
	.S2END(Tile_X13Y9_S2BEGb[7:0]),
	.S4END(Tile_X13Y9_S4BEG[15:0]),
	.SS4END(Tile_X13Y9_SS4BEG[15:0]),
	.W1END(Tile_X14Y10_W1BEG[3:0]),
	.W2MID(Tile_X14Y10_W2BEG[7:0]),
	.W2END(Tile_X14Y10_W2BEGb[7:0]),
	.WW4END(Tile_X14Y10_WW4BEG[15:0]),
	.W6END(Tile_X14Y10_W6BEG[11:0]),
	.N1BEG(Tile_X13Y10_N1BEG[3:0]),
	.N2BEG(Tile_X13Y10_N2BEG[7:0]),
	.N2BEGb(Tile_X13Y10_N2BEGb[7:0]),
	.N4BEG(Tile_X13Y10_N4BEG[15:0]),
	.NN4BEG(Tile_X13Y10_NN4BEG[15:0]),
	.E1BEG(Tile_X13Y10_E1BEG[3:0]),
	.E2BEG(Tile_X13Y10_E2BEG[7:0]),
	.E2BEGb(Tile_X13Y10_E2BEGb[7:0]),
	.EE4BEG(Tile_X13Y10_EE4BEG[15:0]),
	.E6BEG(Tile_X13Y10_E6BEG[11:0]),
	.S1BEG(Tile_X13Y10_S1BEG[3:0]),
	.S2BEG(Tile_X13Y10_S2BEG[7:0]),
	.S2BEGb(Tile_X13Y10_S2BEGb[7:0]),
	.S4BEG(Tile_X13Y10_S4BEG[15:0]),
	.SS4BEG(Tile_X13Y10_SS4BEG[15:0]),
	.W1BEG(Tile_X13Y10_W1BEG[3:0]),
	.W2BEG(Tile_X13Y10_W2BEG[7:0]),
	.W2BEGb(Tile_X13Y10_W2BEGb[7:0]),
	.WW4BEG(Tile_X13Y10_WW4BEG[15:0]),
	.W6BEG(Tile_X13Y10_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X13Y11_UserCLKo),
	.UserCLKo(Tile_X13Y10_UserCLKo),
	.FrameData(Tile_X12Y10_FrameData_O), 
	.FrameData_O(Tile_X13Y10_FrameData_O), 
	.FrameStrobe(Tile_X13Y11_FrameStrobe_O),
	.FrameStrobe_O(Tile_X13Y10_FrameStrobe_O)
	);

	LUT4AB Tile_X14Y10_LUT4AB (
	.N1END(Tile_X14Y11_N1BEG[3:0]),
	.N2MID(Tile_X14Y11_N2BEG[7:0]),
	.N2END(Tile_X14Y11_N2BEGb[7:0]),
	.N4END(Tile_X14Y11_N4BEG[15:0]),
	.NN4END(Tile_X14Y11_NN4BEG[15:0]),
	.Ci(Tile_X14Y11_Co[0:0]),
	.E1END(Tile_X13Y10_E1BEG[3:0]),
	.E2MID(Tile_X13Y10_E2BEG[7:0]),
	.E2END(Tile_X13Y10_E2BEGb[7:0]),
	.EE4END(Tile_X13Y10_EE4BEG[15:0]),
	.E6END(Tile_X13Y10_E6BEG[11:0]),
	.S1END(Tile_X14Y9_S1BEG[3:0]),
	.S2MID(Tile_X14Y9_S2BEG[7:0]),
	.S2END(Tile_X14Y9_S2BEGb[7:0]),
	.S4END(Tile_X14Y9_S4BEG[15:0]),
	.SS4END(Tile_X14Y9_SS4BEG[15:0]),
	.W1END(Tile_X15Y10_W1BEG[3:0]),
	.W2MID(Tile_X15Y10_W2BEG[7:0]),
	.W2END(Tile_X15Y10_W2BEGb[7:0]),
	.WW4END(Tile_X15Y10_WW4BEG[15:0]),
	.W6END(Tile_X15Y10_W6BEG[11:0]),
	.N1BEG(Tile_X14Y10_N1BEG[3:0]),
	.N2BEG(Tile_X14Y10_N2BEG[7:0]),
	.N2BEGb(Tile_X14Y10_N2BEGb[7:0]),
	.N4BEG(Tile_X14Y10_N4BEG[15:0]),
	.NN4BEG(Tile_X14Y10_NN4BEG[15:0]),
	.Co(Tile_X14Y10_Co[0:0]),
	.E1BEG(Tile_X14Y10_E1BEG[3:0]),
	.E2BEG(Tile_X14Y10_E2BEG[7:0]),
	.E2BEGb(Tile_X14Y10_E2BEGb[7:0]),
	.EE4BEG(Tile_X14Y10_EE4BEG[15:0]),
	.E6BEG(Tile_X14Y10_E6BEG[11:0]),
	.S1BEG(Tile_X14Y10_S1BEG[3:0]),
	.S2BEG(Tile_X14Y10_S2BEG[7:0]),
	.S2BEGb(Tile_X14Y10_S2BEGb[7:0]),
	.S4BEG(Tile_X14Y10_S4BEG[15:0]),
	.SS4BEG(Tile_X14Y10_SS4BEG[15:0]),
	.W1BEG(Tile_X14Y10_W1BEG[3:0]),
	.W2BEG(Tile_X14Y10_W2BEG[7:0]),
	.W2BEGb(Tile_X14Y10_W2BEGb[7:0]),
	.WW4BEG(Tile_X14Y10_WW4BEG[15:0]),
	.W6BEG(Tile_X14Y10_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X14Y11_UserCLKo),
	.UserCLKo(Tile_X14Y10_UserCLKo),
	.FrameData(Tile_X13Y10_FrameData_O), 
	.FrameData_O(Tile_X14Y10_FrameData_O), 
	.FrameStrobe(Tile_X14Y11_FrameStrobe_O),
	.FrameStrobe_O(Tile_X14Y10_FrameStrobe_O)
	);

	RAM_IO Tile_X15Y10_RAM_IO (
	.N1END(Tile_X15Y11_N1BEG[3:0]),
	.N2MID(Tile_X15Y11_N2BEG[7:0]),
	.N2END(Tile_X15Y11_N2BEGb[7:0]),
	.N4END(Tile_X15Y11_N4BEG[15:0]),
	.E1END(Tile_X14Y10_E1BEG[3:0]),
	.E2MID(Tile_X14Y10_E2BEG[7:0]),
	.E2END(Tile_X14Y10_E2BEGb[7:0]),
	.EE4END(Tile_X14Y10_EE4BEG[15:0]),
	.E6END(Tile_X14Y10_E6BEG[11:0]),
	.S1END(Tile_X15Y9_S1BEG[3:0]),
	.S2MID(Tile_X15Y9_S2BEG[7:0]),
	.S2END(Tile_X15Y9_S2BEGb[7:0]),
	.S4END(Tile_X15Y9_S4BEG[15:0]),
	.N1BEG(Tile_X15Y10_N1BEG[3:0]),
	.N2BEG(Tile_X15Y10_N2BEG[7:0]),
	.N2BEGb(Tile_X15Y10_N2BEGb[7:0]),
	.N4BEG(Tile_X15Y10_N4BEG[15:0]),
	.S1BEG(Tile_X15Y10_S1BEG[3:0]),
	.S2BEG(Tile_X15Y10_S2BEG[7:0]),
	.S2BEGb(Tile_X15Y10_S2BEGb[7:0]),
	.S4BEG(Tile_X15Y10_S4BEG[15:0]),
	.W1BEG(Tile_X15Y10_W1BEG[3:0]),
	.W2BEG(Tile_X15Y10_W2BEG[7:0]),
	.W2BEGb(Tile_X15Y10_W2BEGb[7:0]),
	.WW4BEG(Tile_X15Y10_WW4BEG[15:0]),
	.W6BEG(Tile_X15Y10_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.RAM2FAB_D0_I0(Tile_X15Y10_RAM2FAB_D0_I0),
	.RAM2FAB_D0_I1(Tile_X15Y10_RAM2FAB_D0_I1),
	.RAM2FAB_D0_I2(Tile_X15Y10_RAM2FAB_D0_I2),
	.RAM2FAB_D0_I3(Tile_X15Y10_RAM2FAB_D0_I3),
	.UserCLK(Tile_X15Y11_UserCLKo),
	.RAM2FAB_D1_I0(Tile_X15Y10_RAM2FAB_D1_I0),
	.RAM2FAB_D1_I1(Tile_X15Y10_RAM2FAB_D1_I1),
	.RAM2FAB_D1_I2(Tile_X15Y10_RAM2FAB_D1_I2),
	.RAM2FAB_D1_I3(Tile_X15Y10_RAM2FAB_D1_I3),
	.RAM2FAB_D2_I0(Tile_X15Y10_RAM2FAB_D2_I0),
	.RAM2FAB_D2_I1(Tile_X15Y10_RAM2FAB_D2_I1),
	.RAM2FAB_D2_I2(Tile_X15Y10_RAM2FAB_D2_I2),
	.RAM2FAB_D2_I3(Tile_X15Y10_RAM2FAB_D2_I3),
	.RAM2FAB_D3_I0(Tile_X15Y10_RAM2FAB_D3_I0),
	.RAM2FAB_D3_I1(Tile_X15Y10_RAM2FAB_D3_I1),
	.RAM2FAB_D3_I2(Tile_X15Y10_RAM2FAB_D3_I2),
	.RAM2FAB_D3_I3(Tile_X15Y10_RAM2FAB_D3_I3),
	.FAB2RAM_D0_O0(Tile_X15Y10_FAB2RAM_D0_O0),
	.FAB2RAM_D0_O1(Tile_X15Y10_FAB2RAM_D0_O1),
	.FAB2RAM_D0_O2(Tile_X15Y10_FAB2RAM_D0_O2),
	.FAB2RAM_D0_O3(Tile_X15Y10_FAB2RAM_D0_O3),
	.FAB2RAM_D1_O0(Tile_X15Y10_FAB2RAM_D1_O0),
	.FAB2RAM_D1_O1(Tile_X15Y10_FAB2RAM_D1_O1),
	.FAB2RAM_D1_O2(Tile_X15Y10_FAB2RAM_D1_O2),
	.FAB2RAM_D1_O3(Tile_X15Y10_FAB2RAM_D1_O3),
	.FAB2RAM_D2_O0(Tile_X15Y10_FAB2RAM_D2_O0),
	.FAB2RAM_D2_O1(Tile_X15Y10_FAB2RAM_D2_O1),
	.FAB2RAM_D2_O2(Tile_X15Y10_FAB2RAM_D2_O2),
	.FAB2RAM_D2_O3(Tile_X15Y10_FAB2RAM_D2_O3),
	.FAB2RAM_D3_O0(Tile_X15Y10_FAB2RAM_D3_O0),
	.FAB2RAM_D3_O1(Tile_X15Y10_FAB2RAM_D3_O1),
	.FAB2RAM_D3_O2(Tile_X15Y10_FAB2RAM_D3_O2),
	.FAB2RAM_D3_O3(Tile_X15Y10_FAB2RAM_D3_O3),
	.FAB2RAM_A0_O0(Tile_X15Y10_FAB2RAM_A0_O0),
	.FAB2RAM_A0_O1(Tile_X15Y10_FAB2RAM_A0_O1),
	.FAB2RAM_A0_O2(Tile_X15Y10_FAB2RAM_A0_O2),
	.FAB2RAM_A0_O3(Tile_X15Y10_FAB2RAM_A0_O3),
	.FAB2RAM_A1_O0(Tile_X15Y10_FAB2RAM_A1_O0),
	.FAB2RAM_A1_O1(Tile_X15Y10_FAB2RAM_A1_O1),
	.FAB2RAM_A1_O2(Tile_X15Y10_FAB2RAM_A1_O2),
	.FAB2RAM_A1_O3(Tile_X15Y10_FAB2RAM_A1_O3),
	.FAB2RAM_C_O0(Tile_X15Y10_FAB2RAM_C_O0),
	.FAB2RAM_C_O1(Tile_X15Y10_FAB2RAM_C_O1),
	.FAB2RAM_C_O2(Tile_X15Y10_FAB2RAM_C_O2),
	.FAB2RAM_C_O3(Tile_X15Y10_FAB2RAM_C_O3),
	.Config_accessC_bit0(Tile_X15Y10_Config_accessC_bit0),
	.Config_accessC_bit1(Tile_X15Y10_Config_accessC_bit1),
	.Config_accessC_bit2(Tile_X15Y10_Config_accessC_bit2),
	.Config_accessC_bit3(Tile_X15Y10_Config_accessC_bit3),
	.UserCLKo(Tile_X15Y10_UserCLKo),
	.FrameData(Tile_X14Y10_FrameData_O), 
	.FrameData_O(Tile_X15Y10_FrameData_O), 
	.FrameStrobe(Tile_X15Y11_FrameStrobe_O),
	.FrameStrobe_O(Tile_X15Y10_FrameStrobe_O)
	);

	W_IO Tile_X0Y11_W_IO (
	.W1END(Tile_X1Y11_W1BEG[3:0]),
	.W2MID(Tile_X1Y11_W2BEG[7:0]),
	.W2END(Tile_X1Y11_W2BEGb[7:0]),
	.WW4END(Tile_X1Y11_WW4BEG[15:0]),
	.W6END(Tile_X1Y11_W6BEG[11:0]),
	.E1BEG(Tile_X0Y11_E1BEG[3:0]),
	.E2BEG(Tile_X0Y11_E2BEG[7:0]),
	.E2BEGb(Tile_X0Y11_E2BEGb[7:0]),
	.EE4BEG(Tile_X0Y11_EE4BEG[15:0]),
	.E6BEG(Tile_X0Y11_E6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.A_I_top(Tile_X0Y11_A_I_top),
	.A_T_top(Tile_X0Y11_A_T_top),
	.A_O_top(Tile_X0Y11_A_O_top),
	.UserCLK(Tile_X0Y12_UserCLKo),
	.B_I_top(Tile_X0Y11_B_I_top),
	.B_T_top(Tile_X0Y11_B_T_top),
	.B_O_top(Tile_X0Y11_B_O_top),
	.A_config_C_bit0(Tile_X0Y11_A_config_C_bit0),
	.A_config_C_bit1(Tile_X0Y11_A_config_C_bit1),
	.A_config_C_bit2(Tile_X0Y11_A_config_C_bit2),
	.A_config_C_bit3(Tile_X0Y11_A_config_C_bit3),
	.B_config_C_bit0(Tile_X0Y11_B_config_C_bit0),
	.B_config_C_bit1(Tile_X0Y11_B_config_C_bit1),
	.B_config_C_bit2(Tile_X0Y11_B_config_C_bit2),
	.B_config_C_bit3(Tile_X0Y11_B_config_C_bit3),
	.UserCLKo(Tile_X0Y11_UserCLKo),
	.FrameData(Tile_Y11_FrameData), 
	.FrameData_O(Tile_X0Y11_FrameData_O), 
	.FrameStrobe(Tile_X0Y12_FrameStrobe_O),
	.FrameStrobe_O(Tile_X0Y11_FrameStrobe_O)
	);

	LUT4AB Tile_X1Y11_LUT4AB (
	.N1END(Tile_X1Y12_N1BEG[3:0]),
	.N2MID(Tile_X1Y12_N2BEG[7:0]),
	.N2END(Tile_X1Y12_N2BEGb[7:0]),
	.N4END(Tile_X1Y12_N4BEG[15:0]),
	.NN4END(Tile_X1Y12_NN4BEG[15:0]),
	.Ci(Tile_X1Y12_Co[0:0]),
	.E1END(Tile_X0Y11_E1BEG[3:0]),
	.E2MID(Tile_X0Y11_E2BEG[7:0]),
	.E2END(Tile_X0Y11_E2BEGb[7:0]),
	.EE4END(Tile_X0Y11_EE4BEG[15:0]),
	.E6END(Tile_X0Y11_E6BEG[11:0]),
	.S1END(Tile_X1Y10_S1BEG[3:0]),
	.S2MID(Tile_X1Y10_S2BEG[7:0]),
	.S2END(Tile_X1Y10_S2BEGb[7:0]),
	.S4END(Tile_X1Y10_S4BEG[15:0]),
	.SS4END(Tile_X1Y10_SS4BEG[15:0]),
	.W1END(Tile_X2Y11_W1BEG[3:0]),
	.W2MID(Tile_X2Y11_W2BEG[7:0]),
	.W2END(Tile_X2Y11_W2BEGb[7:0]),
	.WW4END(Tile_X2Y11_WW4BEG[15:0]),
	.W6END(Tile_X2Y11_W6BEG[11:0]),
	.N1BEG(Tile_X1Y11_N1BEG[3:0]),
	.N2BEG(Tile_X1Y11_N2BEG[7:0]),
	.N2BEGb(Tile_X1Y11_N2BEGb[7:0]),
	.N4BEG(Tile_X1Y11_N4BEG[15:0]),
	.NN4BEG(Tile_X1Y11_NN4BEG[15:0]),
	.Co(Tile_X1Y11_Co[0:0]),
	.E1BEG(Tile_X1Y11_E1BEG[3:0]),
	.E2BEG(Tile_X1Y11_E2BEG[7:0]),
	.E2BEGb(Tile_X1Y11_E2BEGb[7:0]),
	.EE4BEG(Tile_X1Y11_EE4BEG[15:0]),
	.E6BEG(Tile_X1Y11_E6BEG[11:0]),
	.S1BEG(Tile_X1Y11_S1BEG[3:0]),
	.S2BEG(Tile_X1Y11_S2BEG[7:0]),
	.S2BEGb(Tile_X1Y11_S2BEGb[7:0]),
	.S4BEG(Tile_X1Y11_S4BEG[15:0]),
	.SS4BEG(Tile_X1Y11_SS4BEG[15:0]),
	.W1BEG(Tile_X1Y11_W1BEG[3:0]),
	.W2BEG(Tile_X1Y11_W2BEG[7:0]),
	.W2BEGb(Tile_X1Y11_W2BEGb[7:0]),
	.WW4BEG(Tile_X1Y11_WW4BEG[15:0]),
	.W6BEG(Tile_X1Y11_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X1Y12_UserCLKo),
	.UserCLKo(Tile_X1Y11_UserCLKo),
	.FrameData(Tile_X0Y11_FrameData_O), 
	.FrameData_O(Tile_X1Y11_FrameData_O), 
	.FrameStrobe(Tile_X1Y12_FrameStrobe_O),
	.FrameStrobe_O(Tile_X1Y11_FrameStrobe_O)
	);

	RegFile Tile_X2Y11_RegFile (
	.N1END(Tile_X2Y12_N1BEG[3:0]),
	.N2MID(Tile_X2Y12_N2BEG[7:0]),
	.N2END(Tile_X2Y12_N2BEGb[7:0]),
	.N4END(Tile_X2Y12_N4BEG[15:0]),
	.NN4END(Tile_X2Y12_NN4BEG[15:0]),
	.E1END(Tile_X1Y11_E1BEG[3:0]),
	.E2MID(Tile_X1Y11_E2BEG[7:0]),
	.E2END(Tile_X1Y11_E2BEGb[7:0]),
	.EE4END(Tile_X1Y11_EE4BEG[15:0]),
	.E6END(Tile_X1Y11_E6BEG[11:0]),
	.S1END(Tile_X2Y10_S1BEG[3:0]),
	.S2MID(Tile_X2Y10_S2BEG[7:0]),
	.S2END(Tile_X2Y10_S2BEGb[7:0]),
	.S4END(Tile_X2Y10_S4BEG[15:0]),
	.SS4END(Tile_X2Y10_SS4BEG[15:0]),
	.W1END(Tile_X3Y11_W1BEG[3:0]),
	.W2MID(Tile_X3Y11_W2BEG[7:0]),
	.W2END(Tile_X3Y11_W2BEGb[7:0]),
	.WW4END(Tile_X3Y11_WW4BEG[15:0]),
	.W6END(Tile_X3Y11_W6BEG[11:0]),
	.N1BEG(Tile_X2Y11_N1BEG[3:0]),
	.N2BEG(Tile_X2Y11_N2BEG[7:0]),
	.N2BEGb(Tile_X2Y11_N2BEGb[7:0]),
	.N4BEG(Tile_X2Y11_N4BEG[15:0]),
	.NN4BEG(Tile_X2Y11_NN4BEG[15:0]),
	.E1BEG(Tile_X2Y11_E1BEG[3:0]),
	.E2BEG(Tile_X2Y11_E2BEG[7:0]),
	.E2BEGb(Tile_X2Y11_E2BEGb[7:0]),
	.EE4BEG(Tile_X2Y11_EE4BEG[15:0]),
	.E6BEG(Tile_X2Y11_E6BEG[11:0]),
	.S1BEG(Tile_X2Y11_S1BEG[3:0]),
	.S2BEG(Tile_X2Y11_S2BEG[7:0]),
	.S2BEGb(Tile_X2Y11_S2BEGb[7:0]),
	.S4BEG(Tile_X2Y11_S4BEG[15:0]),
	.SS4BEG(Tile_X2Y11_SS4BEG[15:0]),
	.W1BEG(Tile_X2Y11_W1BEG[3:0]),
	.W2BEG(Tile_X2Y11_W2BEG[7:0]),
	.W2BEGb(Tile_X2Y11_W2BEGb[7:0]),
	.WW4BEG(Tile_X2Y11_WW4BEG[15:0]),
	.W6BEG(Tile_X2Y11_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X2Y12_UserCLKo),
	.UserCLKo(Tile_X2Y11_UserCLKo),
	.FrameData(Tile_X1Y11_FrameData_O), 
	.FrameData_O(Tile_X2Y11_FrameData_O), 
	.FrameStrobe(Tile_X2Y12_FrameStrobe_O),
	.FrameStrobe_O(Tile_X2Y11_FrameStrobe_O)
	);

	LUT4AB Tile_X3Y11_LUT4AB (
	.N1END(Tile_X3Y12_N1BEG[3:0]),
	.N2MID(Tile_X3Y12_N2BEG[7:0]),
	.N2END(Tile_X3Y12_N2BEGb[7:0]),
	.N4END(Tile_X3Y12_N4BEG[15:0]),
	.NN4END(Tile_X3Y12_NN4BEG[15:0]),
	.Ci(Tile_X3Y12_Co[0:0]),
	.E1END(Tile_X2Y11_E1BEG[3:0]),
	.E2MID(Tile_X2Y11_E2BEG[7:0]),
	.E2END(Tile_X2Y11_E2BEGb[7:0]),
	.EE4END(Tile_X2Y11_EE4BEG[15:0]),
	.E6END(Tile_X2Y11_E6BEG[11:0]),
	.S1END(Tile_X3Y10_S1BEG[3:0]),
	.S2MID(Tile_X3Y10_S2BEG[7:0]),
	.S2END(Tile_X3Y10_S2BEGb[7:0]),
	.S4END(Tile_X3Y10_S4BEG[15:0]),
	.SS4END(Tile_X3Y10_SS4BEG[15:0]),
	.W1END(Tile_X4Y11_W1BEG[3:0]),
	.W2MID(Tile_X4Y11_W2BEG[7:0]),
	.W2END(Tile_X4Y11_W2BEGb[7:0]),
	.WW4END(Tile_X4Y11_WW4BEG[15:0]),
	.W6END(Tile_X4Y11_W6BEG[11:0]),
	.N1BEG(Tile_X3Y11_N1BEG[3:0]),
	.N2BEG(Tile_X3Y11_N2BEG[7:0]),
	.N2BEGb(Tile_X3Y11_N2BEGb[7:0]),
	.N4BEG(Tile_X3Y11_N4BEG[15:0]),
	.NN4BEG(Tile_X3Y11_NN4BEG[15:0]),
	.Co(Tile_X3Y11_Co[0:0]),
	.E1BEG(Tile_X3Y11_E1BEG[3:0]),
	.E2BEG(Tile_X3Y11_E2BEG[7:0]),
	.E2BEGb(Tile_X3Y11_E2BEGb[7:0]),
	.EE4BEG(Tile_X3Y11_EE4BEG[15:0]),
	.E6BEG(Tile_X3Y11_E6BEG[11:0]),
	.S1BEG(Tile_X3Y11_S1BEG[3:0]),
	.S2BEG(Tile_X3Y11_S2BEG[7:0]),
	.S2BEGb(Tile_X3Y11_S2BEGb[7:0]),
	.S4BEG(Tile_X3Y11_S4BEG[15:0]),
	.SS4BEG(Tile_X3Y11_SS4BEG[15:0]),
	.W1BEG(Tile_X3Y11_W1BEG[3:0]),
	.W2BEG(Tile_X3Y11_W2BEG[7:0]),
	.W2BEGb(Tile_X3Y11_W2BEGb[7:0]),
	.WW4BEG(Tile_X3Y11_WW4BEG[15:0]),
	.W6BEG(Tile_X3Y11_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X3Y12_UserCLKo),
	.UserCLKo(Tile_X3Y11_UserCLKo),
	.FrameData(Tile_X2Y11_FrameData_O), 
	.FrameData_O(Tile_X3Y11_FrameData_O), 
	.FrameStrobe(Tile_X3Y12_FrameStrobe_O),
	.FrameStrobe_O(Tile_X3Y11_FrameStrobe_O)
	);

	LUT4AB Tile_X4Y11_LUT4AB (
	.N1END(Tile_X4Y12_N1BEG[3:0]),
	.N2MID(Tile_X4Y12_N2BEG[7:0]),
	.N2END(Tile_X4Y12_N2BEGb[7:0]),
	.N4END(Tile_X4Y12_N4BEG[15:0]),
	.NN4END(Tile_X4Y12_NN4BEG[15:0]),
	.Ci(Tile_X4Y12_Co[0:0]),
	.E1END(Tile_X3Y11_E1BEG[3:0]),
	.E2MID(Tile_X3Y11_E2BEG[7:0]),
	.E2END(Tile_X3Y11_E2BEGb[7:0]),
	.EE4END(Tile_X3Y11_EE4BEG[15:0]),
	.E6END(Tile_X3Y11_E6BEG[11:0]),
	.S1END(Tile_X4Y10_S1BEG[3:0]),
	.S2MID(Tile_X4Y10_S2BEG[7:0]),
	.S2END(Tile_X4Y10_S2BEGb[7:0]),
	.S4END(Tile_X4Y10_S4BEG[15:0]),
	.SS4END(Tile_X4Y10_SS4BEG[15:0]),
	.W1END(Tile_X5Y11_W1BEG[3:0]),
	.W2MID(Tile_X5Y11_W2BEG[7:0]),
	.W2END(Tile_X5Y11_W2BEGb[7:0]),
	.WW4END(Tile_X5Y11_WW4BEG[15:0]),
	.W6END(Tile_X5Y11_W6BEG[11:0]),
	.N1BEG(Tile_X4Y11_N1BEG[3:0]),
	.N2BEG(Tile_X4Y11_N2BEG[7:0]),
	.N2BEGb(Tile_X4Y11_N2BEGb[7:0]),
	.N4BEG(Tile_X4Y11_N4BEG[15:0]),
	.NN4BEG(Tile_X4Y11_NN4BEG[15:0]),
	.Co(Tile_X4Y11_Co[0:0]),
	.E1BEG(Tile_X4Y11_E1BEG[3:0]),
	.E2BEG(Tile_X4Y11_E2BEG[7:0]),
	.E2BEGb(Tile_X4Y11_E2BEGb[7:0]),
	.EE4BEG(Tile_X4Y11_EE4BEG[15:0]),
	.E6BEG(Tile_X4Y11_E6BEG[11:0]),
	.S1BEG(Tile_X4Y11_S1BEG[3:0]),
	.S2BEG(Tile_X4Y11_S2BEG[7:0]),
	.S2BEGb(Tile_X4Y11_S2BEGb[7:0]),
	.S4BEG(Tile_X4Y11_S4BEG[15:0]),
	.SS4BEG(Tile_X4Y11_SS4BEG[15:0]),
	.W1BEG(Tile_X4Y11_W1BEG[3:0]),
	.W2BEG(Tile_X4Y11_W2BEG[7:0]),
	.W2BEGb(Tile_X4Y11_W2BEGb[7:0]),
	.WW4BEG(Tile_X4Y11_WW4BEG[15:0]),
	.W6BEG(Tile_X4Y11_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X4Y12_UserCLKo),
	.UserCLKo(Tile_X4Y11_UserCLKo),
	.FrameData(Tile_X3Y11_FrameData_O), 
	.FrameData_O(Tile_X4Y11_FrameData_O), 
	.FrameStrobe(Tile_X4Y12_FrameStrobe_O),
	.FrameStrobe_O(Tile_X4Y11_FrameStrobe_O)
	);


	LUT4AB Tile_X6Y11_LUT4AB (
	.N1END(Tile_X6Y12_N1BEG[3:0]),
	.N2MID(Tile_X6Y12_N2BEG[7:0]),
	.N2END(Tile_X6Y12_N2BEGb[7:0]),
	.N4END(Tile_X6Y12_N4BEG[15:0]),
	.NN4END(Tile_X6Y12_NN4BEG[15:0]),
	.Ci(Tile_X6Y12_Co[0:0]),
	.E1END(Tile_X5Y11_E1BEG[3:0]),
	.E2MID(Tile_X5Y11_E2BEG[7:0]),
	.E2END(Tile_X5Y11_E2BEGb[7:0]),
	.EE4END(Tile_X5Y11_EE4BEG[15:0]),
	.E6END(Tile_X5Y11_E6BEG[11:0]),
	.S1END(Tile_X6Y10_S1BEG[3:0]),
	.S2MID(Tile_X6Y10_S2BEG[7:0]),
	.S2END(Tile_X6Y10_S2BEGb[7:0]),
	.S4END(Tile_X6Y10_S4BEG[15:0]),
	.SS4END(Tile_X6Y10_SS4BEG[15:0]),
	.W1END(Tile_X7Y11_W1BEG[3:0]),
	.W2MID(Tile_X7Y11_W2BEG[7:0]),
	.W2END(Tile_X7Y11_W2BEGb[7:0]),
	.WW4END(Tile_X7Y11_WW4BEG[15:0]),
	.W6END(Tile_X7Y11_W6BEG[11:0]),
	.N1BEG(Tile_X6Y11_N1BEG[3:0]),
	.N2BEG(Tile_X6Y11_N2BEG[7:0]),
	.N2BEGb(Tile_X6Y11_N2BEGb[7:0]),
	.N4BEG(Tile_X6Y11_N4BEG[15:0]),
	.NN4BEG(Tile_X6Y11_NN4BEG[15:0]),
	.Co(Tile_X6Y11_Co[0:0]),
	.E1BEG(Tile_X6Y11_E1BEG[3:0]),
	.E2BEG(Tile_X6Y11_E2BEG[7:0]),
	.E2BEGb(Tile_X6Y11_E2BEGb[7:0]),
	.EE4BEG(Tile_X6Y11_EE4BEG[15:0]),
	.E6BEG(Tile_X6Y11_E6BEG[11:0]),
	.S1BEG(Tile_X6Y11_S1BEG[3:0]),
	.S2BEG(Tile_X6Y11_S2BEG[7:0]),
	.S2BEGb(Tile_X6Y11_S2BEGb[7:0]),
	.S4BEG(Tile_X6Y11_S4BEG[15:0]),
	.SS4BEG(Tile_X6Y11_SS4BEG[15:0]),
	.W1BEG(Tile_X6Y11_W1BEG[3:0]),
	.W2BEG(Tile_X6Y11_W2BEG[7:0]),
	.W2BEGb(Tile_X6Y11_W2BEGb[7:0]),
	.WW4BEG(Tile_X6Y11_WW4BEG[15:0]),
	.W6BEG(Tile_X6Y11_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X6Y12_UserCLKo),
	.UserCLKo(Tile_X6Y11_UserCLKo),
	.FrameData(Tile_X5Y11_FrameData_O), 
	.FrameData_O(Tile_X6Y11_FrameData_O), 
	.FrameStrobe(Tile_X6Y12_FrameStrobe_O),
	.FrameStrobe_O(Tile_X6Y11_FrameStrobe_O)
	);

	LUT4AB Tile_X7Y11_LUT4AB (
	.N1END(Tile_X7Y12_N1BEG[3:0]),
	.N2MID(Tile_X7Y12_N2BEG[7:0]),
	.N2END(Tile_X7Y12_N2BEGb[7:0]),
	.N4END(Tile_X7Y12_N4BEG[15:0]),
	.NN4END(Tile_X7Y12_NN4BEG[15:0]),
	.Ci(Tile_X7Y12_Co[0:0]),
	.E1END(Tile_X6Y11_E1BEG[3:0]),
	.E2MID(Tile_X6Y11_E2BEG[7:0]),
	.E2END(Tile_X6Y11_E2BEGb[7:0]),
	.EE4END(Tile_X6Y11_EE4BEG[15:0]),
	.E6END(Tile_X6Y11_E6BEG[11:0]),
	.S1END(Tile_X7Y10_S1BEG[3:0]),
	.S2MID(Tile_X7Y10_S2BEG[7:0]),
	.S2END(Tile_X7Y10_S2BEGb[7:0]),
	.S4END(Tile_X7Y10_S4BEG[15:0]),
	.SS4END(Tile_X7Y10_SS4BEG[15:0]),
	.W1END(Tile_X8Y11_W1BEG[3:0]),
	.W2MID(Tile_X8Y11_W2BEG[7:0]),
	.W2END(Tile_X8Y11_W2BEGb[7:0]),
	.WW4END(Tile_X8Y11_WW4BEG[15:0]),
	.W6END(Tile_X8Y11_W6BEG[11:0]),
	.N1BEG(Tile_X7Y11_N1BEG[3:0]),
	.N2BEG(Tile_X7Y11_N2BEG[7:0]),
	.N2BEGb(Tile_X7Y11_N2BEGb[7:0]),
	.N4BEG(Tile_X7Y11_N4BEG[15:0]),
	.NN4BEG(Tile_X7Y11_NN4BEG[15:0]),
	.Co(Tile_X7Y11_Co[0:0]),
	.E1BEG(Tile_X7Y11_E1BEG[3:0]),
	.E2BEG(Tile_X7Y11_E2BEG[7:0]),
	.E2BEGb(Tile_X7Y11_E2BEGb[7:0]),
	.EE4BEG(Tile_X7Y11_EE4BEG[15:0]),
	.E6BEG(Tile_X7Y11_E6BEG[11:0]),
	.S1BEG(Tile_X7Y11_S1BEG[3:0]),
	.S2BEG(Tile_X7Y11_S2BEG[7:0]),
	.S2BEGb(Tile_X7Y11_S2BEGb[7:0]),
	.S4BEG(Tile_X7Y11_S4BEG[15:0]),
	.SS4BEG(Tile_X7Y11_SS4BEG[15:0]),
	.W1BEG(Tile_X7Y11_W1BEG[3:0]),
	.W2BEG(Tile_X7Y11_W2BEG[7:0]),
	.W2BEGb(Tile_X7Y11_W2BEGb[7:0]),
	.WW4BEG(Tile_X7Y11_WW4BEG[15:0]),
	.W6BEG(Tile_X7Y11_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X7Y12_UserCLKo),
	.UserCLKo(Tile_X7Y11_UserCLKo),
	.FrameData(Tile_X6Y11_FrameData_O), 
	.FrameData_O(Tile_X7Y11_FrameData_O), 
	.FrameStrobe(Tile_X7Y12_FrameStrobe_O),
	.FrameStrobe_O(Tile_X7Y11_FrameStrobe_O)
	);

	LUT4AB Tile_X8Y11_LUT4AB (
	.N1END(Tile_X8Y12_N1BEG[3:0]),
	.N2MID(Tile_X8Y12_N2BEG[7:0]),
	.N2END(Tile_X8Y12_N2BEGb[7:0]),
	.N4END(Tile_X8Y12_N4BEG[15:0]),
	.NN4END(Tile_X8Y12_NN4BEG[15:0]),
	.Ci(Tile_X8Y12_Co[0:0]),
	.E1END(Tile_X7Y11_E1BEG[3:0]),
	.E2MID(Tile_X7Y11_E2BEG[7:0]),
	.E2END(Tile_X7Y11_E2BEGb[7:0]),
	.EE4END(Tile_X7Y11_EE4BEG[15:0]),
	.E6END(Tile_X7Y11_E6BEG[11:0]),
	.S1END(Tile_X8Y10_S1BEG[3:0]),
	.S2MID(Tile_X8Y10_S2BEG[7:0]),
	.S2END(Tile_X8Y10_S2BEGb[7:0]),
	.S4END(Tile_X8Y10_S4BEG[15:0]),
	.SS4END(Tile_X8Y10_SS4BEG[15:0]),
	.W1END(Tile_X9Y11_W1BEG[3:0]),
	.W2MID(Tile_X9Y11_W2BEG[7:0]),
	.W2END(Tile_X9Y11_W2BEGb[7:0]),
	.WW4END(Tile_X9Y11_WW4BEG[15:0]),
	.W6END(Tile_X9Y11_W6BEG[11:0]),
	.N1BEG(Tile_X8Y11_N1BEG[3:0]),
	.N2BEG(Tile_X8Y11_N2BEG[7:0]),
	.N2BEGb(Tile_X8Y11_N2BEGb[7:0]),
	.N4BEG(Tile_X8Y11_N4BEG[15:0]),
	.NN4BEG(Tile_X8Y11_NN4BEG[15:0]),
	.Co(Tile_X8Y11_Co[0:0]),
	.E1BEG(Tile_X8Y11_E1BEG[3:0]),
	.E2BEG(Tile_X8Y11_E2BEG[7:0]),
	.E2BEGb(Tile_X8Y11_E2BEGb[7:0]),
	.EE4BEG(Tile_X8Y11_EE4BEG[15:0]),
	.E6BEG(Tile_X8Y11_E6BEG[11:0]),
	.S1BEG(Tile_X8Y11_S1BEG[3:0]),
	.S2BEG(Tile_X8Y11_S2BEG[7:0]),
	.S2BEGb(Tile_X8Y11_S2BEGb[7:0]),
	.S4BEG(Tile_X8Y11_S4BEG[15:0]),
	.SS4BEG(Tile_X8Y11_SS4BEG[15:0]),
	.W1BEG(Tile_X8Y11_W1BEG[3:0]),
	.W2BEG(Tile_X8Y11_W2BEG[7:0]),
	.W2BEGb(Tile_X8Y11_W2BEGb[7:0]),
	.WW4BEG(Tile_X8Y11_WW4BEG[15:0]),
	.W6BEG(Tile_X8Y11_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X8Y12_UserCLKo),
	.UserCLKo(Tile_X8Y11_UserCLKo),
	.FrameData(Tile_X7Y11_FrameData_O), 
	.FrameData_O(Tile_X8Y11_FrameData_O), 
	.FrameStrobe(Tile_X8Y12_FrameStrobe_O),
	.FrameStrobe_O(Tile_X8Y11_FrameStrobe_O)
	);


	LUT4AB Tile_X10Y11_LUT4AB (
	.N1END(Tile_X10Y12_N1BEG[3:0]),
	.N2MID(Tile_X10Y12_N2BEG[7:0]),
	.N2END(Tile_X10Y12_N2BEGb[7:0]),
	.N4END(Tile_X10Y12_N4BEG[15:0]),
	.NN4END(Tile_X10Y12_NN4BEG[15:0]),
	.Ci(Tile_X10Y12_Co[0:0]),
	.E1END(Tile_X9Y11_E1BEG[3:0]),
	.E2MID(Tile_X9Y11_E2BEG[7:0]),
	.E2END(Tile_X9Y11_E2BEGb[7:0]),
	.EE4END(Tile_X9Y11_EE4BEG[15:0]),
	.E6END(Tile_X9Y11_E6BEG[11:0]),
	.S1END(Tile_X10Y10_S1BEG[3:0]),
	.S2MID(Tile_X10Y10_S2BEG[7:0]),
	.S2END(Tile_X10Y10_S2BEGb[7:0]),
	.S4END(Tile_X10Y10_S4BEG[15:0]),
	.SS4END(Tile_X10Y10_SS4BEG[15:0]),
	.W1END(Tile_X11Y11_W1BEG[3:0]),
	.W2MID(Tile_X11Y11_W2BEG[7:0]),
	.W2END(Tile_X11Y11_W2BEGb[7:0]),
	.WW4END(Tile_X11Y11_WW4BEG[15:0]),
	.W6END(Tile_X11Y11_W6BEG[11:0]),
	.N1BEG(Tile_X10Y11_N1BEG[3:0]),
	.N2BEG(Tile_X10Y11_N2BEG[7:0]),
	.N2BEGb(Tile_X10Y11_N2BEGb[7:0]),
	.N4BEG(Tile_X10Y11_N4BEG[15:0]),
	.NN4BEG(Tile_X10Y11_NN4BEG[15:0]),
	.Co(Tile_X10Y11_Co[0:0]),
	.E1BEG(Tile_X10Y11_E1BEG[3:0]),
	.E2BEG(Tile_X10Y11_E2BEG[7:0]),
	.E2BEGb(Tile_X10Y11_E2BEGb[7:0]),
	.EE4BEG(Tile_X10Y11_EE4BEG[15:0]),
	.E6BEG(Tile_X10Y11_E6BEG[11:0]),
	.S1BEG(Tile_X10Y11_S1BEG[3:0]),
	.S2BEG(Tile_X10Y11_S2BEG[7:0]),
	.S2BEGb(Tile_X10Y11_S2BEGb[7:0]),
	.S4BEG(Tile_X10Y11_S4BEG[15:0]),
	.SS4BEG(Tile_X10Y11_SS4BEG[15:0]),
	.W1BEG(Tile_X10Y11_W1BEG[3:0]),
	.W2BEG(Tile_X10Y11_W2BEG[7:0]),
	.W2BEGb(Tile_X10Y11_W2BEGb[7:0]),
	.WW4BEG(Tile_X10Y11_WW4BEG[15:0]),
	.W6BEG(Tile_X10Y11_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X10Y12_UserCLKo),
	.UserCLKo(Tile_X10Y11_UserCLKo),
	.FrameData(Tile_X9Y11_FrameData_O), 
	.FrameData_O(Tile_X10Y11_FrameData_O), 
	.FrameStrobe(Tile_X10Y12_FrameStrobe_O),
	.FrameStrobe_O(Tile_X10Y11_FrameStrobe_O)
	);

	LUT4AB Tile_X11Y11_LUT4AB (
	.N1END(Tile_X11Y12_N1BEG[3:0]),
	.N2MID(Tile_X11Y12_N2BEG[7:0]),
	.N2END(Tile_X11Y12_N2BEGb[7:0]),
	.N4END(Tile_X11Y12_N4BEG[15:0]),
	.NN4END(Tile_X11Y12_NN4BEG[15:0]),
	.Ci(Tile_X11Y12_Co[0:0]),
	.E1END(Tile_X10Y11_E1BEG[3:0]),
	.E2MID(Tile_X10Y11_E2BEG[7:0]),
	.E2END(Tile_X10Y11_E2BEGb[7:0]),
	.EE4END(Tile_X10Y11_EE4BEG[15:0]),
	.E6END(Tile_X10Y11_E6BEG[11:0]),
	.S1END(Tile_X11Y10_S1BEG[3:0]),
	.S2MID(Tile_X11Y10_S2BEG[7:0]),
	.S2END(Tile_X11Y10_S2BEGb[7:0]),
	.S4END(Tile_X11Y10_S4BEG[15:0]),
	.SS4END(Tile_X11Y10_SS4BEG[15:0]),
	.W1END(Tile_X12Y11_W1BEG[3:0]),
	.W2MID(Tile_X12Y11_W2BEG[7:0]),
	.W2END(Tile_X12Y11_W2BEGb[7:0]),
	.WW4END(Tile_X12Y11_WW4BEG[15:0]),
	.W6END(Tile_X12Y11_W6BEG[11:0]),
	.N1BEG(Tile_X11Y11_N1BEG[3:0]),
	.N2BEG(Tile_X11Y11_N2BEG[7:0]),
	.N2BEGb(Tile_X11Y11_N2BEGb[7:0]),
	.N4BEG(Tile_X11Y11_N4BEG[15:0]),
	.NN4BEG(Tile_X11Y11_NN4BEG[15:0]),
	.Co(Tile_X11Y11_Co[0:0]),
	.E1BEG(Tile_X11Y11_E1BEG[3:0]),
	.E2BEG(Tile_X11Y11_E2BEG[7:0]),
	.E2BEGb(Tile_X11Y11_E2BEGb[7:0]),
	.EE4BEG(Tile_X11Y11_EE4BEG[15:0]),
	.E6BEG(Tile_X11Y11_E6BEG[11:0]),
	.S1BEG(Tile_X11Y11_S1BEG[3:0]),
	.S2BEG(Tile_X11Y11_S2BEG[7:0]),
	.S2BEGb(Tile_X11Y11_S2BEGb[7:0]),
	.S4BEG(Tile_X11Y11_S4BEG[15:0]),
	.SS4BEG(Tile_X11Y11_SS4BEG[15:0]),
	.W1BEG(Tile_X11Y11_W1BEG[3:0]),
	.W2BEG(Tile_X11Y11_W2BEG[7:0]),
	.W2BEGb(Tile_X11Y11_W2BEGb[7:0]),
	.WW4BEG(Tile_X11Y11_WW4BEG[15:0]),
	.W6BEG(Tile_X11Y11_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X11Y12_UserCLKo),
	.UserCLKo(Tile_X11Y11_UserCLKo),
	.FrameData(Tile_X10Y11_FrameData_O), 
	.FrameData_O(Tile_X11Y11_FrameData_O), 
	.FrameStrobe(Tile_X11Y12_FrameStrobe_O),
	.FrameStrobe_O(Tile_X11Y11_FrameStrobe_O)
	);

	LUT4AB Tile_X12Y11_LUT4AB (
	.N1END(Tile_X12Y12_N1BEG[3:0]),
	.N2MID(Tile_X12Y12_N2BEG[7:0]),
	.N2END(Tile_X12Y12_N2BEGb[7:0]),
	.N4END(Tile_X12Y12_N4BEG[15:0]),
	.NN4END(Tile_X12Y12_NN4BEG[15:0]),
	.Ci(Tile_X12Y12_Co[0:0]),
	.E1END(Tile_X11Y11_E1BEG[3:0]),
	.E2MID(Tile_X11Y11_E2BEG[7:0]),
	.E2END(Tile_X11Y11_E2BEGb[7:0]),
	.EE4END(Tile_X11Y11_EE4BEG[15:0]),
	.E6END(Tile_X11Y11_E6BEG[11:0]),
	.S1END(Tile_X12Y10_S1BEG[3:0]),
	.S2MID(Tile_X12Y10_S2BEG[7:0]),
	.S2END(Tile_X12Y10_S2BEGb[7:0]),
	.S4END(Tile_X12Y10_S4BEG[15:0]),
	.SS4END(Tile_X12Y10_SS4BEG[15:0]),
	.W1END(Tile_X13Y11_W1BEG[3:0]),
	.W2MID(Tile_X13Y11_W2BEG[7:0]),
	.W2END(Tile_X13Y11_W2BEGb[7:0]),
	.WW4END(Tile_X13Y11_WW4BEG[15:0]),
	.W6END(Tile_X13Y11_W6BEG[11:0]),
	.N1BEG(Tile_X12Y11_N1BEG[3:0]),
	.N2BEG(Tile_X12Y11_N2BEG[7:0]),
	.N2BEGb(Tile_X12Y11_N2BEGb[7:0]),
	.N4BEG(Tile_X12Y11_N4BEG[15:0]),
	.NN4BEG(Tile_X12Y11_NN4BEG[15:0]),
	.Co(Tile_X12Y11_Co[0:0]),
	.E1BEG(Tile_X12Y11_E1BEG[3:0]),
	.E2BEG(Tile_X12Y11_E2BEG[7:0]),
	.E2BEGb(Tile_X12Y11_E2BEGb[7:0]),
	.EE4BEG(Tile_X12Y11_EE4BEG[15:0]),
	.E6BEG(Tile_X12Y11_E6BEG[11:0]),
	.S1BEG(Tile_X12Y11_S1BEG[3:0]),
	.S2BEG(Tile_X12Y11_S2BEG[7:0]),
	.S2BEGb(Tile_X12Y11_S2BEGb[7:0]),
	.S4BEG(Tile_X12Y11_S4BEG[15:0]),
	.SS4BEG(Tile_X12Y11_SS4BEG[15:0]),
	.W1BEG(Tile_X12Y11_W1BEG[3:0]),
	.W2BEG(Tile_X12Y11_W2BEG[7:0]),
	.W2BEGb(Tile_X12Y11_W2BEGb[7:0]),
	.WW4BEG(Tile_X12Y11_WW4BEG[15:0]),
	.W6BEG(Tile_X12Y11_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X12Y12_UserCLKo),
	.UserCLKo(Tile_X12Y11_UserCLKo),
	.FrameData(Tile_X11Y11_FrameData_O), 
	.FrameData_O(Tile_X12Y11_FrameData_O), 
	.FrameStrobe(Tile_X12Y12_FrameStrobe_O),
	.FrameStrobe_O(Tile_X12Y11_FrameStrobe_O)
	);

	RegFile Tile_X13Y11_RegFile (
	.N1END(Tile_X13Y12_N1BEG[3:0]),
	.N2MID(Tile_X13Y12_N2BEG[7:0]),
	.N2END(Tile_X13Y12_N2BEGb[7:0]),
	.N4END(Tile_X13Y12_N4BEG[15:0]),
	.NN4END(Tile_X13Y12_NN4BEG[15:0]),
	.E1END(Tile_X12Y11_E1BEG[3:0]),
	.E2MID(Tile_X12Y11_E2BEG[7:0]),
	.E2END(Tile_X12Y11_E2BEGb[7:0]),
	.EE4END(Tile_X12Y11_EE4BEG[15:0]),
	.E6END(Tile_X12Y11_E6BEG[11:0]),
	.S1END(Tile_X13Y10_S1BEG[3:0]),
	.S2MID(Tile_X13Y10_S2BEG[7:0]),
	.S2END(Tile_X13Y10_S2BEGb[7:0]),
	.S4END(Tile_X13Y10_S4BEG[15:0]),
	.SS4END(Tile_X13Y10_SS4BEG[15:0]),
	.W1END(Tile_X14Y11_W1BEG[3:0]),
	.W2MID(Tile_X14Y11_W2BEG[7:0]),
	.W2END(Tile_X14Y11_W2BEGb[7:0]),
	.WW4END(Tile_X14Y11_WW4BEG[15:0]),
	.W6END(Tile_X14Y11_W6BEG[11:0]),
	.N1BEG(Tile_X13Y11_N1BEG[3:0]),
	.N2BEG(Tile_X13Y11_N2BEG[7:0]),
	.N2BEGb(Tile_X13Y11_N2BEGb[7:0]),
	.N4BEG(Tile_X13Y11_N4BEG[15:0]),
	.NN4BEG(Tile_X13Y11_NN4BEG[15:0]),
	.E1BEG(Tile_X13Y11_E1BEG[3:0]),
	.E2BEG(Tile_X13Y11_E2BEG[7:0]),
	.E2BEGb(Tile_X13Y11_E2BEGb[7:0]),
	.EE4BEG(Tile_X13Y11_EE4BEG[15:0]),
	.E6BEG(Tile_X13Y11_E6BEG[11:0]),
	.S1BEG(Tile_X13Y11_S1BEG[3:0]),
	.S2BEG(Tile_X13Y11_S2BEG[7:0]),
	.S2BEGb(Tile_X13Y11_S2BEGb[7:0]),
	.S4BEG(Tile_X13Y11_S4BEG[15:0]),
	.SS4BEG(Tile_X13Y11_SS4BEG[15:0]),
	.W1BEG(Tile_X13Y11_W1BEG[3:0]),
	.W2BEG(Tile_X13Y11_W2BEG[7:0]),
	.W2BEGb(Tile_X13Y11_W2BEGb[7:0]),
	.WW4BEG(Tile_X13Y11_WW4BEG[15:0]),
	.W6BEG(Tile_X13Y11_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X13Y12_UserCLKo),
	.UserCLKo(Tile_X13Y11_UserCLKo),
	.FrameData(Tile_X12Y11_FrameData_O), 
	.FrameData_O(Tile_X13Y11_FrameData_O), 
	.FrameStrobe(Tile_X13Y12_FrameStrobe_O),
	.FrameStrobe_O(Tile_X13Y11_FrameStrobe_O)
	);

	LUT4AB Tile_X14Y11_LUT4AB (
	.N1END(Tile_X14Y12_N1BEG[3:0]),
	.N2MID(Tile_X14Y12_N2BEG[7:0]),
	.N2END(Tile_X14Y12_N2BEGb[7:0]),
	.N4END(Tile_X14Y12_N4BEG[15:0]),
	.NN4END(Tile_X14Y12_NN4BEG[15:0]),
	.Ci(Tile_X14Y12_Co[0:0]),
	.E1END(Tile_X13Y11_E1BEG[3:0]),
	.E2MID(Tile_X13Y11_E2BEG[7:0]),
	.E2END(Tile_X13Y11_E2BEGb[7:0]),
	.EE4END(Tile_X13Y11_EE4BEG[15:0]),
	.E6END(Tile_X13Y11_E6BEG[11:0]),
	.S1END(Tile_X14Y10_S1BEG[3:0]),
	.S2MID(Tile_X14Y10_S2BEG[7:0]),
	.S2END(Tile_X14Y10_S2BEGb[7:0]),
	.S4END(Tile_X14Y10_S4BEG[15:0]),
	.SS4END(Tile_X14Y10_SS4BEG[15:0]),
	.W1END(Tile_X15Y11_W1BEG[3:0]),
	.W2MID(Tile_X15Y11_W2BEG[7:0]),
	.W2END(Tile_X15Y11_W2BEGb[7:0]),
	.WW4END(Tile_X15Y11_WW4BEG[15:0]),
	.W6END(Tile_X15Y11_W6BEG[11:0]),
	.N1BEG(Tile_X14Y11_N1BEG[3:0]),
	.N2BEG(Tile_X14Y11_N2BEG[7:0]),
	.N2BEGb(Tile_X14Y11_N2BEGb[7:0]),
	.N4BEG(Tile_X14Y11_N4BEG[15:0]),
	.NN4BEG(Tile_X14Y11_NN4BEG[15:0]),
	.Co(Tile_X14Y11_Co[0:0]),
	.E1BEG(Tile_X14Y11_E1BEG[3:0]),
	.E2BEG(Tile_X14Y11_E2BEG[7:0]),
	.E2BEGb(Tile_X14Y11_E2BEGb[7:0]),
	.EE4BEG(Tile_X14Y11_EE4BEG[15:0]),
	.E6BEG(Tile_X14Y11_E6BEG[11:0]),
	.S1BEG(Tile_X14Y11_S1BEG[3:0]),
	.S2BEG(Tile_X14Y11_S2BEG[7:0]),
	.S2BEGb(Tile_X14Y11_S2BEGb[7:0]),
	.S4BEG(Tile_X14Y11_S4BEG[15:0]),
	.SS4BEG(Tile_X14Y11_SS4BEG[15:0]),
	.W1BEG(Tile_X14Y11_W1BEG[3:0]),
	.W2BEG(Tile_X14Y11_W2BEG[7:0]),
	.W2BEGb(Tile_X14Y11_W2BEGb[7:0]),
	.WW4BEG(Tile_X14Y11_WW4BEG[15:0]),
	.W6BEG(Tile_X14Y11_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X14Y12_UserCLKo),
	.UserCLKo(Tile_X14Y11_UserCLKo),
	.FrameData(Tile_X13Y11_FrameData_O), 
	.FrameData_O(Tile_X14Y11_FrameData_O), 
	.FrameStrobe(Tile_X14Y12_FrameStrobe_O),
	.FrameStrobe_O(Tile_X14Y11_FrameStrobe_O)
	);

	RAM_IO Tile_X15Y11_RAM_IO (
	.N1END(Tile_X15Y12_N1BEG[3:0]),
	.N2MID(Tile_X15Y12_N2BEG[7:0]),
	.N2END(Tile_X15Y12_N2BEGb[7:0]),
	.N4END(Tile_X15Y12_N4BEG[15:0]),
	.E1END(Tile_X14Y11_E1BEG[3:0]),
	.E2MID(Tile_X14Y11_E2BEG[7:0]),
	.E2END(Tile_X14Y11_E2BEGb[7:0]),
	.EE4END(Tile_X14Y11_EE4BEG[15:0]),
	.E6END(Tile_X14Y11_E6BEG[11:0]),
	.S1END(Tile_X15Y10_S1BEG[3:0]),
	.S2MID(Tile_X15Y10_S2BEG[7:0]),
	.S2END(Tile_X15Y10_S2BEGb[7:0]),
	.S4END(Tile_X15Y10_S4BEG[15:0]),
	.N1BEG(Tile_X15Y11_N1BEG[3:0]),
	.N2BEG(Tile_X15Y11_N2BEG[7:0]),
	.N2BEGb(Tile_X15Y11_N2BEGb[7:0]),
	.N4BEG(Tile_X15Y11_N4BEG[15:0]),
	.S1BEG(Tile_X15Y11_S1BEG[3:0]),
	.S2BEG(Tile_X15Y11_S2BEG[7:0]),
	.S2BEGb(Tile_X15Y11_S2BEGb[7:0]),
	.S4BEG(Tile_X15Y11_S4BEG[15:0]),
	.W1BEG(Tile_X15Y11_W1BEG[3:0]),
	.W2BEG(Tile_X15Y11_W2BEG[7:0]),
	.W2BEGb(Tile_X15Y11_W2BEGb[7:0]),
	.WW4BEG(Tile_X15Y11_WW4BEG[15:0]),
	.W6BEG(Tile_X15Y11_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.RAM2FAB_D0_I0(Tile_X15Y11_RAM2FAB_D0_I0),
	.RAM2FAB_D0_I1(Tile_X15Y11_RAM2FAB_D0_I1),
	.RAM2FAB_D0_I2(Tile_X15Y11_RAM2FAB_D0_I2),
	.RAM2FAB_D0_I3(Tile_X15Y11_RAM2FAB_D0_I3),
	.UserCLK(Tile_X15Y12_UserCLKo),
	.RAM2FAB_D1_I0(Tile_X15Y11_RAM2FAB_D1_I0),
	.RAM2FAB_D1_I1(Tile_X15Y11_RAM2FAB_D1_I1),
	.RAM2FAB_D1_I2(Tile_X15Y11_RAM2FAB_D1_I2),
	.RAM2FAB_D1_I3(Tile_X15Y11_RAM2FAB_D1_I3),
	.RAM2FAB_D2_I0(Tile_X15Y11_RAM2FAB_D2_I0),
	.RAM2FAB_D2_I1(Tile_X15Y11_RAM2FAB_D2_I1),
	.RAM2FAB_D2_I2(Tile_X15Y11_RAM2FAB_D2_I2),
	.RAM2FAB_D2_I3(Tile_X15Y11_RAM2FAB_D2_I3),
	.RAM2FAB_D3_I0(Tile_X15Y11_RAM2FAB_D3_I0),
	.RAM2FAB_D3_I1(Tile_X15Y11_RAM2FAB_D3_I1),
	.RAM2FAB_D3_I2(Tile_X15Y11_RAM2FAB_D3_I2),
	.RAM2FAB_D3_I3(Tile_X15Y11_RAM2FAB_D3_I3),
	.FAB2RAM_D0_O0(Tile_X15Y11_FAB2RAM_D0_O0),
	.FAB2RAM_D0_O1(Tile_X15Y11_FAB2RAM_D0_O1),
	.FAB2RAM_D0_O2(Tile_X15Y11_FAB2RAM_D0_O2),
	.FAB2RAM_D0_O3(Tile_X15Y11_FAB2RAM_D0_O3),
	.FAB2RAM_D1_O0(Tile_X15Y11_FAB2RAM_D1_O0),
	.FAB2RAM_D1_O1(Tile_X15Y11_FAB2RAM_D1_O1),
	.FAB2RAM_D1_O2(Tile_X15Y11_FAB2RAM_D1_O2),
	.FAB2RAM_D1_O3(Tile_X15Y11_FAB2RAM_D1_O3),
	.FAB2RAM_D2_O0(Tile_X15Y11_FAB2RAM_D2_O0),
	.FAB2RAM_D2_O1(Tile_X15Y11_FAB2RAM_D2_O1),
	.FAB2RAM_D2_O2(Tile_X15Y11_FAB2RAM_D2_O2),
	.FAB2RAM_D2_O3(Tile_X15Y11_FAB2RAM_D2_O3),
	.FAB2RAM_D3_O0(Tile_X15Y11_FAB2RAM_D3_O0),
	.FAB2RAM_D3_O1(Tile_X15Y11_FAB2RAM_D3_O1),
	.FAB2RAM_D3_O2(Tile_X15Y11_FAB2RAM_D3_O2),
	.FAB2RAM_D3_O3(Tile_X15Y11_FAB2RAM_D3_O3),
	.FAB2RAM_A0_O0(Tile_X15Y11_FAB2RAM_A0_O0),
	.FAB2RAM_A0_O1(Tile_X15Y11_FAB2RAM_A0_O1),
	.FAB2RAM_A0_O2(Tile_X15Y11_FAB2RAM_A0_O2),
	.FAB2RAM_A0_O3(Tile_X15Y11_FAB2RAM_A0_O3),
	.FAB2RAM_A1_O0(Tile_X15Y11_FAB2RAM_A1_O0),
	.FAB2RAM_A1_O1(Tile_X15Y11_FAB2RAM_A1_O1),
	.FAB2RAM_A1_O2(Tile_X15Y11_FAB2RAM_A1_O2),
	.FAB2RAM_A1_O3(Tile_X15Y11_FAB2RAM_A1_O3),
	.FAB2RAM_C_O0(Tile_X15Y11_FAB2RAM_C_O0),
	.FAB2RAM_C_O1(Tile_X15Y11_FAB2RAM_C_O1),
	.FAB2RAM_C_O2(Tile_X15Y11_FAB2RAM_C_O2),
	.FAB2RAM_C_O3(Tile_X15Y11_FAB2RAM_C_O3),
	.Config_accessC_bit0(Tile_X15Y11_Config_accessC_bit0),
	.Config_accessC_bit1(Tile_X15Y11_Config_accessC_bit1),
	.Config_accessC_bit2(Tile_X15Y11_Config_accessC_bit2),
	.Config_accessC_bit3(Tile_X15Y11_Config_accessC_bit3),
	.UserCLKo(Tile_X15Y11_UserCLKo),
	.FrameData(Tile_X14Y11_FrameData_O), 
	.FrameData_O(Tile_X15Y11_FrameData_O), 
	.FrameStrobe(Tile_X15Y12_FrameStrobe_O),
	.FrameStrobe_O(Tile_X15Y11_FrameStrobe_O)
	);

	W_IO Tile_X0Y12_W_IO (
	.W1END(Tile_X1Y12_W1BEG[3:0]),
	.W2MID(Tile_X1Y12_W2BEG[7:0]),
	.W2END(Tile_X1Y12_W2BEGb[7:0]),
	.WW4END(Tile_X1Y12_WW4BEG[15:0]),
	.W6END(Tile_X1Y12_W6BEG[11:0]),
	.E1BEG(Tile_X0Y12_E1BEG[3:0]),
	.E2BEG(Tile_X0Y12_E2BEG[7:0]),
	.E2BEGb(Tile_X0Y12_E2BEGb[7:0]),
	.EE4BEG(Tile_X0Y12_EE4BEG[15:0]),
	.E6BEG(Tile_X0Y12_E6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.A_I_top(Tile_X0Y12_A_I_top),
	.A_T_top(Tile_X0Y12_A_T_top),
	.A_O_top(Tile_X0Y12_A_O_top),
	.UserCLK(UserCLK),
	.B_I_top(Tile_X0Y12_B_I_top),
	.B_T_top(Tile_X0Y12_B_T_top),
	.B_O_top(Tile_X0Y12_B_O_top),
	.A_config_C_bit0(Tile_X0Y12_A_config_C_bit0),
	.A_config_C_bit1(Tile_X0Y12_A_config_C_bit1),
	.A_config_C_bit2(Tile_X0Y12_A_config_C_bit2),
	.A_config_C_bit3(Tile_X0Y12_A_config_C_bit3),
	.B_config_C_bit0(Tile_X0Y12_B_config_C_bit0),
	.B_config_C_bit1(Tile_X0Y12_B_config_C_bit1),
	.B_config_C_bit2(Tile_X0Y12_B_config_C_bit2),
	.B_config_C_bit3(Tile_X0Y12_B_config_C_bit3),
	.UserCLKo(Tile_X0Y12_UserCLKo),
	.FrameData(Tile_Y12_FrameData), 
	.FrameData_O(Tile_X0Y12_FrameData_O), 
	.FrameStrobe(Tile_X0_FrameStrobe),
	.FrameStrobe_O(Tile_X0Y12_FrameStrobe_O)
	);

	LUT4AB Tile_X1Y12_LUT4AB (
	.N1END(Tile_X1Y13_N1BEG[3:0]),
	.N2MID(Tile_X1Y13_N2BEG[7:0]),
	.N2END(Tile_X1Y13_N2BEGb[7:0]),
	.N4END(Tile_X1Y13_N4BEG[15:0]),
	.NN4END(Tile_X1Y13_NN4BEG[15:0]),
	.Ci(Tile_X1Y13_Co[0:0]),
	.E1END(Tile_X0Y12_E1BEG[3:0]),
	.E2MID(Tile_X0Y12_E2BEG[7:0]),
	.E2END(Tile_X0Y12_E2BEGb[7:0]),
	.EE4END(Tile_X0Y12_EE4BEG[15:0]),
	.E6END(Tile_X0Y12_E6BEG[11:0]),
	.S1END(Tile_X1Y11_S1BEG[3:0]),
	.S2MID(Tile_X1Y11_S2BEG[7:0]),
	.S2END(Tile_X1Y11_S2BEGb[7:0]),
	.S4END(Tile_X1Y11_S4BEG[15:0]),
	.SS4END(Tile_X1Y11_SS4BEG[15:0]),
	.W1END(Tile_X2Y12_W1BEG[3:0]),
	.W2MID(Tile_X2Y12_W2BEG[7:0]),
	.W2END(Tile_X2Y12_W2BEGb[7:0]),
	.WW4END(Tile_X2Y12_WW4BEG[15:0]),
	.W6END(Tile_X2Y12_W6BEG[11:0]),
	.N1BEG(Tile_X1Y12_N1BEG[3:0]),
	.N2BEG(Tile_X1Y12_N2BEG[7:0]),
	.N2BEGb(Tile_X1Y12_N2BEGb[7:0]),
	.N4BEG(Tile_X1Y12_N4BEG[15:0]),
	.NN4BEG(Tile_X1Y12_NN4BEG[15:0]),
	.Co(Tile_X1Y12_Co[0:0]),
	.E1BEG(Tile_X1Y12_E1BEG[3:0]),
	.E2BEG(Tile_X1Y12_E2BEG[7:0]),
	.E2BEGb(Tile_X1Y12_E2BEGb[7:0]),
	.EE4BEG(Tile_X1Y12_EE4BEG[15:0]),
	.E6BEG(Tile_X1Y12_E6BEG[11:0]),
	.S1BEG(Tile_X1Y12_S1BEG[3:0]),
	.S2BEG(Tile_X1Y12_S2BEG[7:0]),
	.S2BEGb(Tile_X1Y12_S2BEGb[7:0]),
	.S4BEG(Tile_X1Y12_S4BEG[15:0]),
	.SS4BEG(Tile_X1Y12_SS4BEG[15:0]),
	.W1BEG(Tile_X1Y12_W1BEG[3:0]),
	.W2BEG(Tile_X1Y12_W2BEG[7:0]),
	.W2BEGb(Tile_X1Y12_W2BEGb[7:0]),
	.WW4BEG(Tile_X1Y12_WW4BEG[15:0]),
	.W6BEG(Tile_X1Y12_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X1Y13_UserCLKo),
	.UserCLKo(Tile_X1Y12_UserCLKo),
	.FrameData(Tile_X0Y12_FrameData_O), 
	.FrameData_O(Tile_X1Y12_FrameData_O), 
	.FrameStrobe(Tile_X1Y13_FrameStrobe_O),
	.FrameStrobe_O(Tile_X1Y12_FrameStrobe_O)
	);

	RegFile Tile_X2Y12_RegFile (
	.N1END(Tile_X2Y13_N1BEG[3:0]),
	.N2MID(Tile_X2Y13_N2BEG[7:0]),
	.N2END(Tile_X2Y13_N2BEGb[7:0]),
	.N4END(Tile_X2Y13_N4BEG[15:0]),
	.NN4END(Tile_X2Y13_NN4BEG[15:0]),
	.E1END(Tile_X1Y12_E1BEG[3:0]),
	.E2MID(Tile_X1Y12_E2BEG[7:0]),
	.E2END(Tile_X1Y12_E2BEGb[7:0]),
	.EE4END(Tile_X1Y12_EE4BEG[15:0]),
	.E6END(Tile_X1Y12_E6BEG[11:0]),
	.S1END(Tile_X2Y11_S1BEG[3:0]),
	.S2MID(Tile_X2Y11_S2BEG[7:0]),
	.S2END(Tile_X2Y11_S2BEGb[7:0]),
	.S4END(Tile_X2Y11_S4BEG[15:0]),
	.SS4END(Tile_X2Y11_SS4BEG[15:0]),
	.W1END(Tile_X3Y12_W1BEG[3:0]),
	.W2MID(Tile_X3Y12_W2BEG[7:0]),
	.W2END(Tile_X3Y12_W2BEGb[7:0]),
	.WW4END(Tile_X3Y12_WW4BEG[15:0]),
	.W6END(Tile_X3Y12_W6BEG[11:0]),
	.N1BEG(Tile_X2Y12_N1BEG[3:0]),
	.N2BEG(Tile_X2Y12_N2BEG[7:0]),
	.N2BEGb(Tile_X2Y12_N2BEGb[7:0]),
	.N4BEG(Tile_X2Y12_N4BEG[15:0]),
	.NN4BEG(Tile_X2Y12_NN4BEG[15:0]),
	.E1BEG(Tile_X2Y12_E1BEG[3:0]),
	.E2BEG(Tile_X2Y12_E2BEG[7:0]),
	.E2BEGb(Tile_X2Y12_E2BEGb[7:0]),
	.EE4BEG(Tile_X2Y12_EE4BEG[15:0]),
	.E6BEG(Tile_X2Y12_E6BEG[11:0]),
	.S1BEG(Tile_X2Y12_S1BEG[3:0]),
	.S2BEG(Tile_X2Y12_S2BEG[7:0]),
	.S2BEGb(Tile_X2Y12_S2BEGb[7:0]),
	.S4BEG(Tile_X2Y12_S4BEG[15:0]),
	.SS4BEG(Tile_X2Y12_SS4BEG[15:0]),
	.W1BEG(Tile_X2Y12_W1BEG[3:0]),
	.W2BEG(Tile_X2Y12_W2BEG[7:0]),
	.W2BEGb(Tile_X2Y12_W2BEGb[7:0]),
	.WW4BEG(Tile_X2Y12_WW4BEG[15:0]),
	.W6BEG(Tile_X2Y12_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X2Y13_UserCLKo),
	.UserCLKo(Tile_X2Y12_UserCLKo),
	.FrameData(Tile_X1Y12_FrameData_O), 
	.FrameData_O(Tile_X2Y12_FrameData_O), 
	.FrameStrobe(Tile_X2Y13_FrameStrobe_O),
	.FrameStrobe_O(Tile_X2Y12_FrameStrobe_O)
	);

	LUT4AB Tile_X3Y12_LUT4AB (
	.N1END(Tile_X3Y13_N1BEG[3:0]),
	.N2MID(Tile_X3Y13_N2BEG[7:0]),
	.N2END(Tile_X3Y13_N2BEGb[7:0]),
	.N4END(Tile_X3Y13_N4BEG[15:0]),
	.NN4END(Tile_X3Y13_NN4BEG[15:0]),
	.Ci(Tile_X3Y13_Co[0:0]),
	.E1END(Tile_X2Y12_E1BEG[3:0]),
	.E2MID(Tile_X2Y12_E2BEG[7:0]),
	.E2END(Tile_X2Y12_E2BEGb[7:0]),
	.EE4END(Tile_X2Y12_EE4BEG[15:0]),
	.E6END(Tile_X2Y12_E6BEG[11:0]),
	.S1END(Tile_X3Y11_S1BEG[3:0]),
	.S2MID(Tile_X3Y11_S2BEG[7:0]),
	.S2END(Tile_X3Y11_S2BEGb[7:0]),
	.S4END(Tile_X3Y11_S4BEG[15:0]),
	.SS4END(Tile_X3Y11_SS4BEG[15:0]),
	.W1END(Tile_X4Y12_W1BEG[3:0]),
	.W2MID(Tile_X4Y12_W2BEG[7:0]),
	.W2END(Tile_X4Y12_W2BEGb[7:0]),
	.WW4END(Tile_X4Y12_WW4BEG[15:0]),
	.W6END(Tile_X4Y12_W6BEG[11:0]),
	.N1BEG(Tile_X3Y12_N1BEG[3:0]),
	.N2BEG(Tile_X3Y12_N2BEG[7:0]),
	.N2BEGb(Tile_X3Y12_N2BEGb[7:0]),
	.N4BEG(Tile_X3Y12_N4BEG[15:0]),
	.NN4BEG(Tile_X3Y12_NN4BEG[15:0]),
	.Co(Tile_X3Y12_Co[0:0]),
	.E1BEG(Tile_X3Y12_E1BEG[3:0]),
	.E2BEG(Tile_X3Y12_E2BEG[7:0]),
	.E2BEGb(Tile_X3Y12_E2BEGb[7:0]),
	.EE4BEG(Tile_X3Y12_EE4BEG[15:0]),
	.E6BEG(Tile_X3Y12_E6BEG[11:0]),
	.S1BEG(Tile_X3Y12_S1BEG[3:0]),
	.S2BEG(Tile_X3Y12_S2BEG[7:0]),
	.S2BEGb(Tile_X3Y12_S2BEGb[7:0]),
	.S4BEG(Tile_X3Y12_S4BEG[15:0]),
	.SS4BEG(Tile_X3Y12_SS4BEG[15:0]),
	.W1BEG(Tile_X3Y12_W1BEG[3:0]),
	.W2BEG(Tile_X3Y12_W2BEG[7:0]),
	.W2BEGb(Tile_X3Y12_W2BEGb[7:0]),
	.WW4BEG(Tile_X3Y12_WW4BEG[15:0]),
	.W6BEG(Tile_X3Y12_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X3Y13_UserCLKo),
	.UserCLKo(Tile_X3Y12_UserCLKo),
	.FrameData(Tile_X2Y12_FrameData_O), 
	.FrameData_O(Tile_X3Y12_FrameData_O), 
	.FrameStrobe(Tile_X3Y13_FrameStrobe_O),
	.FrameStrobe_O(Tile_X3Y12_FrameStrobe_O)
	);

	LUT4AB Tile_X4Y12_LUT4AB (
	.N1END(Tile_X4Y13_N1BEG[3:0]),
	.N2MID(Tile_X4Y13_N2BEG[7:0]),
	.N2END(Tile_X4Y13_N2BEGb[7:0]),
	.N4END(Tile_X4Y13_N4BEG[15:0]),
	.NN4END(Tile_X4Y13_NN4BEG[15:0]),
	.Ci(Tile_X4Y13_Co[0:0]),
	.E1END(Tile_X3Y12_E1BEG[3:0]),
	.E2MID(Tile_X3Y12_E2BEG[7:0]),
	.E2END(Tile_X3Y12_E2BEGb[7:0]),
	.EE4END(Tile_X3Y12_EE4BEG[15:0]),
	.E6END(Tile_X3Y12_E6BEG[11:0]),
	.S1END(Tile_X4Y11_S1BEG[3:0]),
	.S2MID(Tile_X4Y11_S2BEG[7:0]),
	.S2END(Tile_X4Y11_S2BEGb[7:0]),
	.S4END(Tile_X4Y11_S4BEG[15:0]),
	.SS4END(Tile_X4Y11_SS4BEG[15:0]),
	.W1END(Tile_X5Y12_W1BEG[3:0]),
	.W2MID(Tile_X5Y12_W2BEG[7:0]),
	.W2END(Tile_X5Y12_W2BEGb[7:0]),
	.WW4END(Tile_X5Y12_WW4BEG[15:0]),
	.W6END(Tile_X5Y12_W6BEG[11:0]),
	.N1BEG(Tile_X4Y12_N1BEG[3:0]),
	.N2BEG(Tile_X4Y12_N2BEG[7:0]),
	.N2BEGb(Tile_X4Y12_N2BEGb[7:0]),
	.N4BEG(Tile_X4Y12_N4BEG[15:0]),
	.NN4BEG(Tile_X4Y12_NN4BEG[15:0]),
	.Co(Tile_X4Y12_Co[0:0]),
	.E1BEG(Tile_X4Y12_E1BEG[3:0]),
	.E2BEG(Tile_X4Y12_E2BEG[7:0]),
	.E2BEGb(Tile_X4Y12_E2BEGb[7:0]),
	.EE4BEG(Tile_X4Y12_EE4BEG[15:0]),
	.E6BEG(Tile_X4Y12_E6BEG[11:0]),
	.S1BEG(Tile_X4Y12_S1BEG[3:0]),
	.S2BEG(Tile_X4Y12_S2BEG[7:0]),
	.S2BEGb(Tile_X4Y12_S2BEGb[7:0]),
	.S4BEG(Tile_X4Y12_S4BEG[15:0]),
	.SS4BEG(Tile_X4Y12_SS4BEG[15:0]),
	.W1BEG(Tile_X4Y12_W1BEG[3:0]),
	.W2BEG(Tile_X4Y12_W2BEG[7:0]),
	.W2BEGb(Tile_X4Y12_W2BEGb[7:0]),
	.WW4BEG(Tile_X4Y12_WW4BEG[15:0]),
	.W6BEG(Tile_X4Y12_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X4Y13_UserCLKo),
	.UserCLKo(Tile_X4Y12_UserCLKo),
	.FrameData(Tile_X3Y12_FrameData_O), 
	.FrameData_O(Tile_X4Y12_FrameData_O), 
	.FrameStrobe(Tile_X4Y13_FrameStrobe_O),
	.FrameStrobe_O(Tile_X4Y12_FrameStrobe_O)
	);


	LUT4AB Tile_X6Y12_LUT4AB (
	.N1END(Tile_X6Y13_N1BEG[3:0]),
	.N2MID(Tile_X6Y13_N2BEG[7:0]),
	.N2END(Tile_X6Y13_N2BEGb[7:0]),
	.N4END(Tile_X6Y13_N4BEG[15:0]),
	.NN4END(Tile_X6Y13_NN4BEG[15:0]),
	.Ci(Tile_X6Y13_Co[0:0]),
	.E1END(Tile_X5Y12_E1BEG[3:0]),
	.E2MID(Tile_X5Y12_E2BEG[7:0]),
	.E2END(Tile_X5Y12_E2BEGb[7:0]),
	.EE4END(Tile_X5Y12_EE4BEG[15:0]),
	.E6END(Tile_X5Y12_E6BEG[11:0]),
	.S1END(Tile_X6Y11_S1BEG[3:0]),
	.S2MID(Tile_X6Y11_S2BEG[7:0]),
	.S2END(Tile_X6Y11_S2BEGb[7:0]),
	.S4END(Tile_X6Y11_S4BEG[15:0]),
	.SS4END(Tile_X6Y11_SS4BEG[15:0]),
	.W1END(Tile_X7Y12_W1BEG[3:0]),
	.W2MID(Tile_X7Y12_W2BEG[7:0]),
	.W2END(Tile_X7Y12_W2BEGb[7:0]),
	.WW4END(Tile_X7Y12_WW4BEG[15:0]),
	.W6END(Tile_X7Y12_W6BEG[11:0]),
	.N1BEG(Tile_X6Y12_N1BEG[3:0]),
	.N2BEG(Tile_X6Y12_N2BEG[7:0]),
	.N2BEGb(Tile_X6Y12_N2BEGb[7:0]),
	.N4BEG(Tile_X6Y12_N4BEG[15:0]),
	.NN4BEG(Tile_X6Y12_NN4BEG[15:0]),
	.Co(Tile_X6Y12_Co[0:0]),
	.E1BEG(Tile_X6Y12_E1BEG[3:0]),
	.E2BEG(Tile_X6Y12_E2BEG[7:0]),
	.E2BEGb(Tile_X6Y12_E2BEGb[7:0]),
	.EE4BEG(Tile_X6Y12_EE4BEG[15:0]),
	.E6BEG(Tile_X6Y12_E6BEG[11:0]),
	.S1BEG(Tile_X6Y12_S1BEG[3:0]),
	.S2BEG(Tile_X6Y12_S2BEG[7:0]),
	.S2BEGb(Tile_X6Y12_S2BEGb[7:0]),
	.S4BEG(Tile_X6Y12_S4BEG[15:0]),
	.SS4BEG(Tile_X6Y12_SS4BEG[15:0]),
	.W1BEG(Tile_X6Y12_W1BEG[3:0]),
	.W2BEG(Tile_X6Y12_W2BEG[7:0]),
	.W2BEGb(Tile_X6Y12_W2BEGb[7:0]),
	.WW4BEG(Tile_X6Y12_WW4BEG[15:0]),
	.W6BEG(Tile_X6Y12_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X6Y13_UserCLKo),
	.UserCLKo(Tile_X6Y12_UserCLKo),
	.FrameData(Tile_X5Y12_FrameData_O), 
	.FrameData_O(Tile_X6Y12_FrameData_O), 
	.FrameStrobe(Tile_X6Y13_FrameStrobe_O),
	.FrameStrobe_O(Tile_X6Y12_FrameStrobe_O)
	);

	LUT4AB Tile_X7Y12_LUT4AB (
	.N1END(Tile_X7Y13_N1BEG[3:0]),
	.N2MID(Tile_X7Y13_N2BEG[7:0]),
	.N2END(Tile_X7Y13_N2BEGb[7:0]),
	.N4END(Tile_X7Y13_N4BEG[15:0]),
	.NN4END(Tile_X7Y13_NN4BEG[15:0]),
	.Ci(Tile_X7Y13_Co[0:0]),
	.E1END(Tile_X6Y12_E1BEG[3:0]),
	.E2MID(Tile_X6Y12_E2BEG[7:0]),
	.E2END(Tile_X6Y12_E2BEGb[7:0]),
	.EE4END(Tile_X6Y12_EE4BEG[15:0]),
	.E6END(Tile_X6Y12_E6BEG[11:0]),
	.S1END(Tile_X7Y11_S1BEG[3:0]),
	.S2MID(Tile_X7Y11_S2BEG[7:0]),
	.S2END(Tile_X7Y11_S2BEGb[7:0]),
	.S4END(Tile_X7Y11_S4BEG[15:0]),
	.SS4END(Tile_X7Y11_SS4BEG[15:0]),
	.W1END(Tile_X8Y12_W1BEG[3:0]),
	.W2MID(Tile_X8Y12_W2BEG[7:0]),
	.W2END(Tile_X8Y12_W2BEGb[7:0]),
	.WW4END(Tile_X8Y12_WW4BEG[15:0]),
	.W6END(Tile_X8Y12_W6BEG[11:0]),
	.N1BEG(Tile_X7Y12_N1BEG[3:0]),
	.N2BEG(Tile_X7Y12_N2BEG[7:0]),
	.N2BEGb(Tile_X7Y12_N2BEGb[7:0]),
	.N4BEG(Tile_X7Y12_N4BEG[15:0]),
	.NN4BEG(Tile_X7Y12_NN4BEG[15:0]),
	.Co(Tile_X7Y12_Co[0:0]),
	.E1BEG(Tile_X7Y12_E1BEG[3:0]),
	.E2BEG(Tile_X7Y12_E2BEG[7:0]),
	.E2BEGb(Tile_X7Y12_E2BEGb[7:0]),
	.EE4BEG(Tile_X7Y12_EE4BEG[15:0]),
	.E6BEG(Tile_X7Y12_E6BEG[11:0]),
	.S1BEG(Tile_X7Y12_S1BEG[3:0]),
	.S2BEG(Tile_X7Y12_S2BEG[7:0]),
	.S2BEGb(Tile_X7Y12_S2BEGb[7:0]),
	.S4BEG(Tile_X7Y12_S4BEG[15:0]),
	.SS4BEG(Tile_X7Y12_SS4BEG[15:0]),
	.W1BEG(Tile_X7Y12_W1BEG[3:0]),
	.W2BEG(Tile_X7Y12_W2BEG[7:0]),
	.W2BEGb(Tile_X7Y12_W2BEGb[7:0]),
	.WW4BEG(Tile_X7Y12_WW4BEG[15:0]),
	.W6BEG(Tile_X7Y12_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X7Y13_UserCLKo),
	.UserCLKo(Tile_X7Y12_UserCLKo),
	.FrameData(Tile_X6Y12_FrameData_O), 
	.FrameData_O(Tile_X7Y12_FrameData_O), 
	.FrameStrobe(Tile_X7Y13_FrameStrobe_O),
	.FrameStrobe_O(Tile_X7Y12_FrameStrobe_O)
	);

	LUT4AB Tile_X8Y12_LUT4AB (
	.N1END(Tile_X8Y13_N1BEG[3:0]),
	.N2MID(Tile_X8Y13_N2BEG[7:0]),
	.N2END(Tile_X8Y13_N2BEGb[7:0]),
	.N4END(Tile_X8Y13_N4BEG[15:0]),
	.NN4END(Tile_X8Y13_NN4BEG[15:0]),
	.Ci(Tile_X8Y13_Co[0:0]),
	.E1END(Tile_X7Y12_E1BEG[3:0]),
	.E2MID(Tile_X7Y12_E2BEG[7:0]),
	.E2END(Tile_X7Y12_E2BEGb[7:0]),
	.EE4END(Tile_X7Y12_EE4BEG[15:0]),
	.E6END(Tile_X7Y12_E6BEG[11:0]),
	.S1END(Tile_X8Y11_S1BEG[3:0]),
	.S2MID(Tile_X8Y11_S2BEG[7:0]),
	.S2END(Tile_X8Y11_S2BEGb[7:0]),
	.S4END(Tile_X8Y11_S4BEG[15:0]),
	.SS4END(Tile_X8Y11_SS4BEG[15:0]),
	.W1END(Tile_X9Y12_W1BEG[3:0]),
	.W2MID(Tile_X9Y12_W2BEG[7:0]),
	.W2END(Tile_X9Y12_W2BEGb[7:0]),
	.WW4END(Tile_X9Y12_WW4BEG[15:0]),
	.W6END(Tile_X9Y12_W6BEG[11:0]),
	.N1BEG(Tile_X8Y12_N1BEG[3:0]),
	.N2BEG(Tile_X8Y12_N2BEG[7:0]),
	.N2BEGb(Tile_X8Y12_N2BEGb[7:0]),
	.N4BEG(Tile_X8Y12_N4BEG[15:0]),
	.NN4BEG(Tile_X8Y12_NN4BEG[15:0]),
	.Co(Tile_X8Y12_Co[0:0]),
	.E1BEG(Tile_X8Y12_E1BEG[3:0]),
	.E2BEG(Tile_X8Y12_E2BEG[7:0]),
	.E2BEGb(Tile_X8Y12_E2BEGb[7:0]),
	.EE4BEG(Tile_X8Y12_EE4BEG[15:0]),
	.E6BEG(Tile_X8Y12_E6BEG[11:0]),
	.S1BEG(Tile_X8Y12_S1BEG[3:0]),
	.S2BEG(Tile_X8Y12_S2BEG[7:0]),
	.S2BEGb(Tile_X8Y12_S2BEGb[7:0]),
	.S4BEG(Tile_X8Y12_S4BEG[15:0]),
	.SS4BEG(Tile_X8Y12_SS4BEG[15:0]),
	.W1BEG(Tile_X8Y12_W1BEG[3:0]),
	.W2BEG(Tile_X8Y12_W2BEG[7:0]),
	.W2BEGb(Tile_X8Y12_W2BEGb[7:0]),
	.WW4BEG(Tile_X8Y12_WW4BEG[15:0]),
	.W6BEG(Tile_X8Y12_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X8Y13_UserCLKo),
	.UserCLKo(Tile_X8Y12_UserCLKo),
	.FrameData(Tile_X7Y12_FrameData_O), 
	.FrameData_O(Tile_X8Y12_FrameData_O), 
	.FrameStrobe(Tile_X8Y13_FrameStrobe_O),
	.FrameStrobe_O(Tile_X8Y12_FrameStrobe_O)
	);


	LUT4AB Tile_X10Y12_LUT4AB (
	.N1END(Tile_X10Y13_N1BEG[3:0]),
	.N2MID(Tile_X10Y13_N2BEG[7:0]),
	.N2END(Tile_X10Y13_N2BEGb[7:0]),
	.N4END(Tile_X10Y13_N4BEG[15:0]),
	.NN4END(Tile_X10Y13_NN4BEG[15:0]),
	.Ci(Tile_X10Y13_Co[0:0]),
	.E1END(Tile_X9Y12_E1BEG[3:0]),
	.E2MID(Tile_X9Y12_E2BEG[7:0]),
	.E2END(Tile_X9Y12_E2BEGb[7:0]),
	.EE4END(Tile_X9Y12_EE4BEG[15:0]),
	.E6END(Tile_X9Y12_E6BEG[11:0]),
	.S1END(Tile_X10Y11_S1BEG[3:0]),
	.S2MID(Tile_X10Y11_S2BEG[7:0]),
	.S2END(Tile_X10Y11_S2BEGb[7:0]),
	.S4END(Tile_X10Y11_S4BEG[15:0]),
	.SS4END(Tile_X10Y11_SS4BEG[15:0]),
	.W1END(Tile_X11Y12_W1BEG[3:0]),
	.W2MID(Tile_X11Y12_W2BEG[7:0]),
	.W2END(Tile_X11Y12_W2BEGb[7:0]),
	.WW4END(Tile_X11Y12_WW4BEG[15:0]),
	.W6END(Tile_X11Y12_W6BEG[11:0]),
	.N1BEG(Tile_X10Y12_N1BEG[3:0]),
	.N2BEG(Tile_X10Y12_N2BEG[7:0]),
	.N2BEGb(Tile_X10Y12_N2BEGb[7:0]),
	.N4BEG(Tile_X10Y12_N4BEG[15:0]),
	.NN4BEG(Tile_X10Y12_NN4BEG[15:0]),
	.Co(Tile_X10Y12_Co[0:0]),
	.E1BEG(Tile_X10Y12_E1BEG[3:0]),
	.E2BEG(Tile_X10Y12_E2BEG[7:0]),
	.E2BEGb(Tile_X10Y12_E2BEGb[7:0]),
	.EE4BEG(Tile_X10Y12_EE4BEG[15:0]),
	.E6BEG(Tile_X10Y12_E6BEG[11:0]),
	.S1BEG(Tile_X10Y12_S1BEG[3:0]),
	.S2BEG(Tile_X10Y12_S2BEG[7:0]),
	.S2BEGb(Tile_X10Y12_S2BEGb[7:0]),
	.S4BEG(Tile_X10Y12_S4BEG[15:0]),
	.SS4BEG(Tile_X10Y12_SS4BEG[15:0]),
	.W1BEG(Tile_X10Y12_W1BEG[3:0]),
	.W2BEG(Tile_X10Y12_W2BEG[7:0]),
	.W2BEGb(Tile_X10Y12_W2BEGb[7:0]),
	.WW4BEG(Tile_X10Y12_WW4BEG[15:0]),
	.W6BEG(Tile_X10Y12_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X10Y13_UserCLKo),
	.UserCLKo(Tile_X10Y12_UserCLKo),
	.FrameData(Tile_X9Y12_FrameData_O), 
	.FrameData_O(Tile_X10Y12_FrameData_O), 
	.FrameStrobe(Tile_X10Y13_FrameStrobe_O),
	.FrameStrobe_O(Tile_X10Y12_FrameStrobe_O)
	);

	LUT4AB Tile_X11Y12_LUT4AB (
	.N1END(Tile_X11Y13_N1BEG[3:0]),
	.N2MID(Tile_X11Y13_N2BEG[7:0]),
	.N2END(Tile_X11Y13_N2BEGb[7:0]),
	.N4END(Tile_X11Y13_N4BEG[15:0]),
	.NN4END(Tile_X11Y13_NN4BEG[15:0]),
	.Ci(Tile_X11Y13_Co[0:0]),
	.E1END(Tile_X10Y12_E1BEG[3:0]),
	.E2MID(Tile_X10Y12_E2BEG[7:0]),
	.E2END(Tile_X10Y12_E2BEGb[7:0]),
	.EE4END(Tile_X10Y12_EE4BEG[15:0]),
	.E6END(Tile_X10Y12_E6BEG[11:0]),
	.S1END(Tile_X11Y11_S1BEG[3:0]),
	.S2MID(Tile_X11Y11_S2BEG[7:0]),
	.S2END(Tile_X11Y11_S2BEGb[7:0]),
	.S4END(Tile_X11Y11_S4BEG[15:0]),
	.SS4END(Tile_X11Y11_SS4BEG[15:0]),
	.W1END(Tile_X12Y12_W1BEG[3:0]),
	.W2MID(Tile_X12Y12_W2BEG[7:0]),
	.W2END(Tile_X12Y12_W2BEGb[7:0]),
	.WW4END(Tile_X12Y12_WW4BEG[15:0]),
	.W6END(Tile_X12Y12_W6BEG[11:0]),
	.N1BEG(Tile_X11Y12_N1BEG[3:0]),
	.N2BEG(Tile_X11Y12_N2BEG[7:0]),
	.N2BEGb(Tile_X11Y12_N2BEGb[7:0]),
	.N4BEG(Tile_X11Y12_N4BEG[15:0]),
	.NN4BEG(Tile_X11Y12_NN4BEG[15:0]),
	.Co(Tile_X11Y12_Co[0:0]),
	.E1BEG(Tile_X11Y12_E1BEG[3:0]),
	.E2BEG(Tile_X11Y12_E2BEG[7:0]),
	.E2BEGb(Tile_X11Y12_E2BEGb[7:0]),
	.EE4BEG(Tile_X11Y12_EE4BEG[15:0]),
	.E6BEG(Tile_X11Y12_E6BEG[11:0]),
	.S1BEG(Tile_X11Y12_S1BEG[3:0]),
	.S2BEG(Tile_X11Y12_S2BEG[7:0]),
	.S2BEGb(Tile_X11Y12_S2BEGb[7:0]),
	.S4BEG(Tile_X11Y12_S4BEG[15:0]),
	.SS4BEG(Tile_X11Y12_SS4BEG[15:0]),
	.W1BEG(Tile_X11Y12_W1BEG[3:0]),
	.W2BEG(Tile_X11Y12_W2BEG[7:0]),
	.W2BEGb(Tile_X11Y12_W2BEGb[7:0]),
	.WW4BEG(Tile_X11Y12_WW4BEG[15:0]),
	.W6BEG(Tile_X11Y12_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X11Y13_UserCLKo),
	.UserCLKo(Tile_X11Y12_UserCLKo),
	.FrameData(Tile_X10Y12_FrameData_O), 
	.FrameData_O(Tile_X11Y12_FrameData_O), 
	.FrameStrobe(Tile_X11Y13_FrameStrobe_O),
	.FrameStrobe_O(Tile_X11Y12_FrameStrobe_O)
	);

	LUT4AB Tile_X12Y12_LUT4AB (
	.N1END(Tile_X12Y13_N1BEG[3:0]),
	.N2MID(Tile_X12Y13_N2BEG[7:0]),
	.N2END(Tile_X12Y13_N2BEGb[7:0]),
	.N4END(Tile_X12Y13_N4BEG[15:0]),
	.NN4END(Tile_X12Y13_NN4BEG[15:0]),
	.Ci(Tile_X12Y13_Co[0:0]),
	.E1END(Tile_X11Y12_E1BEG[3:0]),
	.E2MID(Tile_X11Y12_E2BEG[7:0]),
	.E2END(Tile_X11Y12_E2BEGb[7:0]),
	.EE4END(Tile_X11Y12_EE4BEG[15:0]),
	.E6END(Tile_X11Y12_E6BEG[11:0]),
	.S1END(Tile_X12Y11_S1BEG[3:0]),
	.S2MID(Tile_X12Y11_S2BEG[7:0]),
	.S2END(Tile_X12Y11_S2BEGb[7:0]),
	.S4END(Tile_X12Y11_S4BEG[15:0]),
	.SS4END(Tile_X12Y11_SS4BEG[15:0]),
	.W1END(Tile_X13Y12_W1BEG[3:0]),
	.W2MID(Tile_X13Y12_W2BEG[7:0]),
	.W2END(Tile_X13Y12_W2BEGb[7:0]),
	.WW4END(Tile_X13Y12_WW4BEG[15:0]),
	.W6END(Tile_X13Y12_W6BEG[11:0]),
	.N1BEG(Tile_X12Y12_N1BEG[3:0]),
	.N2BEG(Tile_X12Y12_N2BEG[7:0]),
	.N2BEGb(Tile_X12Y12_N2BEGb[7:0]),
	.N4BEG(Tile_X12Y12_N4BEG[15:0]),
	.NN4BEG(Tile_X12Y12_NN4BEG[15:0]),
	.Co(Tile_X12Y12_Co[0:0]),
	.E1BEG(Tile_X12Y12_E1BEG[3:0]),
	.E2BEG(Tile_X12Y12_E2BEG[7:0]),
	.E2BEGb(Tile_X12Y12_E2BEGb[7:0]),
	.EE4BEG(Tile_X12Y12_EE4BEG[15:0]),
	.E6BEG(Tile_X12Y12_E6BEG[11:0]),
	.S1BEG(Tile_X12Y12_S1BEG[3:0]),
	.S2BEG(Tile_X12Y12_S2BEG[7:0]),
	.S2BEGb(Tile_X12Y12_S2BEGb[7:0]),
	.S4BEG(Tile_X12Y12_S4BEG[15:0]),
	.SS4BEG(Tile_X12Y12_SS4BEG[15:0]),
	.W1BEG(Tile_X12Y12_W1BEG[3:0]),
	.W2BEG(Tile_X12Y12_W2BEG[7:0]),
	.W2BEGb(Tile_X12Y12_W2BEGb[7:0]),
	.WW4BEG(Tile_X12Y12_WW4BEG[15:0]),
	.W6BEG(Tile_X12Y12_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X12Y13_UserCLKo),
	.UserCLKo(Tile_X12Y12_UserCLKo),
	.FrameData(Tile_X11Y12_FrameData_O), 
	.FrameData_O(Tile_X12Y12_FrameData_O), 
	.FrameStrobe(Tile_X12Y13_FrameStrobe_O),
	.FrameStrobe_O(Tile_X12Y12_FrameStrobe_O)
	);

	RegFile Tile_X13Y12_RegFile (
	.N1END(Tile_X13Y13_N1BEG[3:0]),
	.N2MID(Tile_X13Y13_N2BEG[7:0]),
	.N2END(Tile_X13Y13_N2BEGb[7:0]),
	.N4END(Tile_X13Y13_N4BEG[15:0]),
	.NN4END(Tile_X13Y13_NN4BEG[15:0]),
	.E1END(Tile_X12Y12_E1BEG[3:0]),
	.E2MID(Tile_X12Y12_E2BEG[7:0]),
	.E2END(Tile_X12Y12_E2BEGb[7:0]),
	.EE4END(Tile_X12Y12_EE4BEG[15:0]),
	.E6END(Tile_X12Y12_E6BEG[11:0]),
	.S1END(Tile_X13Y11_S1BEG[3:0]),
	.S2MID(Tile_X13Y11_S2BEG[7:0]),
	.S2END(Tile_X13Y11_S2BEGb[7:0]),
	.S4END(Tile_X13Y11_S4BEG[15:0]),
	.SS4END(Tile_X13Y11_SS4BEG[15:0]),
	.W1END(Tile_X14Y12_W1BEG[3:0]),
	.W2MID(Tile_X14Y12_W2BEG[7:0]),
	.W2END(Tile_X14Y12_W2BEGb[7:0]),
	.WW4END(Tile_X14Y12_WW4BEG[15:0]),
	.W6END(Tile_X14Y12_W6BEG[11:0]),
	.N1BEG(Tile_X13Y12_N1BEG[3:0]),
	.N2BEG(Tile_X13Y12_N2BEG[7:0]),
	.N2BEGb(Tile_X13Y12_N2BEGb[7:0]),
	.N4BEG(Tile_X13Y12_N4BEG[15:0]),
	.NN4BEG(Tile_X13Y12_NN4BEG[15:0]),
	.E1BEG(Tile_X13Y12_E1BEG[3:0]),
	.E2BEG(Tile_X13Y12_E2BEG[7:0]),
	.E2BEGb(Tile_X13Y12_E2BEGb[7:0]),
	.EE4BEG(Tile_X13Y12_EE4BEG[15:0]),
	.E6BEG(Tile_X13Y12_E6BEG[11:0]),
	.S1BEG(Tile_X13Y12_S1BEG[3:0]),
	.S2BEG(Tile_X13Y12_S2BEG[7:0]),
	.S2BEGb(Tile_X13Y12_S2BEGb[7:0]),
	.S4BEG(Tile_X13Y12_S4BEG[15:0]),
	.SS4BEG(Tile_X13Y12_SS4BEG[15:0]),
	.W1BEG(Tile_X13Y12_W1BEG[3:0]),
	.W2BEG(Tile_X13Y12_W2BEG[7:0]),
	.W2BEGb(Tile_X13Y12_W2BEGb[7:0]),
	.WW4BEG(Tile_X13Y12_WW4BEG[15:0]),
	.W6BEG(Tile_X13Y12_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X13Y13_UserCLKo),
	.UserCLKo(Tile_X13Y12_UserCLKo),
	.FrameData(Tile_X12Y12_FrameData_O), 
	.FrameData_O(Tile_X13Y12_FrameData_O), 
	.FrameStrobe(Tile_X13Y13_FrameStrobe_O),
	.FrameStrobe_O(Tile_X13Y12_FrameStrobe_O)
	);

	LUT4AB Tile_X14Y12_LUT4AB (
	.N1END(Tile_X14Y13_N1BEG[3:0]),
	.N2MID(Tile_X14Y13_N2BEG[7:0]),
	.N2END(Tile_X14Y13_N2BEGb[7:0]),
	.N4END(Tile_X14Y13_N4BEG[15:0]),
	.NN4END(Tile_X14Y13_NN4BEG[15:0]),
	.Ci(Tile_X14Y13_Co[0:0]),
	.E1END(Tile_X13Y12_E1BEG[3:0]),
	.E2MID(Tile_X13Y12_E2BEG[7:0]),
	.E2END(Tile_X13Y12_E2BEGb[7:0]),
	.EE4END(Tile_X13Y12_EE4BEG[15:0]),
	.E6END(Tile_X13Y12_E6BEG[11:0]),
	.S1END(Tile_X14Y11_S1BEG[3:0]),
	.S2MID(Tile_X14Y11_S2BEG[7:0]),
	.S2END(Tile_X14Y11_S2BEGb[7:0]),
	.S4END(Tile_X14Y11_S4BEG[15:0]),
	.SS4END(Tile_X14Y11_SS4BEG[15:0]),
	.W1END(Tile_X15Y12_W1BEG[3:0]),
	.W2MID(Tile_X15Y12_W2BEG[7:0]),
	.W2END(Tile_X15Y12_W2BEGb[7:0]),
	.WW4END(Tile_X15Y12_WW4BEG[15:0]),
	.W6END(Tile_X15Y12_W6BEG[11:0]),
	.N1BEG(Tile_X14Y12_N1BEG[3:0]),
	.N2BEG(Tile_X14Y12_N2BEG[7:0]),
	.N2BEGb(Tile_X14Y12_N2BEGb[7:0]),
	.N4BEG(Tile_X14Y12_N4BEG[15:0]),
	.NN4BEG(Tile_X14Y12_NN4BEG[15:0]),
	.Co(Tile_X14Y12_Co[0:0]),
	.E1BEG(Tile_X14Y12_E1BEG[3:0]),
	.E2BEG(Tile_X14Y12_E2BEG[7:0]),
	.E2BEGb(Tile_X14Y12_E2BEGb[7:0]),
	.EE4BEG(Tile_X14Y12_EE4BEG[15:0]),
	.E6BEG(Tile_X14Y12_E6BEG[11:0]),
	.S1BEG(Tile_X14Y12_S1BEG[3:0]),
	.S2BEG(Tile_X14Y12_S2BEG[7:0]),
	.S2BEGb(Tile_X14Y12_S2BEGb[7:0]),
	.S4BEG(Tile_X14Y12_S4BEG[15:0]),
	.SS4BEG(Tile_X14Y12_SS4BEG[15:0]),
	.W1BEG(Tile_X14Y12_W1BEG[3:0]),
	.W2BEG(Tile_X14Y12_W2BEG[7:0]),
	.W2BEGb(Tile_X14Y12_W2BEGb[7:0]),
	.WW4BEG(Tile_X14Y12_WW4BEG[15:0]),
	.W6BEG(Tile_X14Y12_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(Tile_X14Y13_UserCLKo),
	.UserCLKo(Tile_X14Y12_UserCLKo),
	.FrameData(Tile_X13Y12_FrameData_O), 
	.FrameData_O(Tile_X14Y12_FrameData_O), 
	.FrameStrobe(Tile_X14Y13_FrameStrobe_O),
	.FrameStrobe_O(Tile_X14Y12_FrameStrobe_O)
	);

	RAM_IO Tile_X15Y12_RAM_IO (
	.N1END(Tile_X15Y13_N1BEG[3:0]),
	.N2MID(Tile_X15Y13_N2BEG[7:0]),
	.N2END(Tile_X15Y13_N2BEGb[7:0]),
	.N4END(Tile_X15Y13_N4BEG[15:0]),
	.E1END(Tile_X14Y12_E1BEG[3:0]),
	.E2MID(Tile_X14Y12_E2BEG[7:0]),
	.E2END(Tile_X14Y12_E2BEGb[7:0]),
	.EE4END(Tile_X14Y12_EE4BEG[15:0]),
	.E6END(Tile_X14Y12_E6BEG[11:0]),
	.S1END(Tile_X15Y11_S1BEG[3:0]),
	.S2MID(Tile_X15Y11_S2BEG[7:0]),
	.S2END(Tile_X15Y11_S2BEGb[7:0]),
	.S4END(Tile_X15Y11_S4BEG[15:0]),
	.N1BEG(Tile_X15Y12_N1BEG[3:0]),
	.N2BEG(Tile_X15Y12_N2BEG[7:0]),
	.N2BEGb(Tile_X15Y12_N2BEGb[7:0]),
	.N4BEG(Tile_X15Y12_N4BEG[15:0]),
	.S1BEG(Tile_X15Y12_S1BEG[3:0]),
	.S2BEG(Tile_X15Y12_S2BEG[7:0]),
	.S2BEGb(Tile_X15Y12_S2BEGb[7:0]),
	.S4BEG(Tile_X15Y12_S4BEG[15:0]),
	.W1BEG(Tile_X15Y12_W1BEG[3:0]),
	.W2BEG(Tile_X15Y12_W2BEG[7:0]),
	.W2BEGb(Tile_X15Y12_W2BEGb[7:0]),
	.WW4BEG(Tile_X15Y12_WW4BEG[15:0]),
	.W6BEG(Tile_X15Y12_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.RAM2FAB_D0_I0(Tile_X15Y12_RAM2FAB_D0_I0),
	.RAM2FAB_D0_I1(Tile_X15Y12_RAM2FAB_D0_I1),
	.RAM2FAB_D0_I2(Tile_X15Y12_RAM2FAB_D0_I2),
	.RAM2FAB_D0_I3(Tile_X15Y12_RAM2FAB_D0_I3),
	.UserCLK(Tile_X15Y13_UserCLKo),
	.RAM2FAB_D1_I0(Tile_X15Y12_RAM2FAB_D1_I0),
	.RAM2FAB_D1_I1(Tile_X15Y12_RAM2FAB_D1_I1),
	.RAM2FAB_D1_I2(Tile_X15Y12_RAM2FAB_D1_I2),
	.RAM2FAB_D1_I3(Tile_X15Y12_RAM2FAB_D1_I3),
	.RAM2FAB_D2_I0(Tile_X15Y12_RAM2FAB_D2_I0),
	.RAM2FAB_D2_I1(Tile_X15Y12_RAM2FAB_D2_I1),
	.RAM2FAB_D2_I2(Tile_X15Y12_RAM2FAB_D2_I2),
	.RAM2FAB_D2_I3(Tile_X15Y12_RAM2FAB_D2_I3),
	.RAM2FAB_D3_I0(Tile_X15Y12_RAM2FAB_D3_I0),
	.RAM2FAB_D3_I1(Tile_X15Y12_RAM2FAB_D3_I1),
	.RAM2FAB_D3_I2(Tile_X15Y12_RAM2FAB_D3_I2),
	.RAM2FAB_D3_I3(Tile_X15Y12_RAM2FAB_D3_I3),
	.FAB2RAM_D0_O0(Tile_X15Y12_FAB2RAM_D0_O0),
	.FAB2RAM_D0_O1(Tile_X15Y12_FAB2RAM_D0_O1),
	.FAB2RAM_D0_O2(Tile_X15Y12_FAB2RAM_D0_O2),
	.FAB2RAM_D0_O3(Tile_X15Y12_FAB2RAM_D0_O3),
	.FAB2RAM_D1_O0(Tile_X15Y12_FAB2RAM_D1_O0),
	.FAB2RAM_D1_O1(Tile_X15Y12_FAB2RAM_D1_O1),
	.FAB2RAM_D1_O2(Tile_X15Y12_FAB2RAM_D1_O2),
	.FAB2RAM_D1_O3(Tile_X15Y12_FAB2RAM_D1_O3),
	.FAB2RAM_D2_O0(Tile_X15Y12_FAB2RAM_D2_O0),
	.FAB2RAM_D2_O1(Tile_X15Y12_FAB2RAM_D2_O1),
	.FAB2RAM_D2_O2(Tile_X15Y12_FAB2RAM_D2_O2),
	.FAB2RAM_D2_O3(Tile_X15Y12_FAB2RAM_D2_O3),
	.FAB2RAM_D3_O0(Tile_X15Y12_FAB2RAM_D3_O0),
	.FAB2RAM_D3_O1(Tile_X15Y12_FAB2RAM_D3_O1),
	.FAB2RAM_D3_O2(Tile_X15Y12_FAB2RAM_D3_O2),
	.FAB2RAM_D3_O3(Tile_X15Y12_FAB2RAM_D3_O3),
	.FAB2RAM_A0_O0(Tile_X15Y12_FAB2RAM_A0_O0),
	.FAB2RAM_A0_O1(Tile_X15Y12_FAB2RAM_A0_O1),
	.FAB2RAM_A0_O2(Tile_X15Y12_FAB2RAM_A0_O2),
	.FAB2RAM_A0_O3(Tile_X15Y12_FAB2RAM_A0_O3),
	.FAB2RAM_A1_O0(Tile_X15Y12_FAB2RAM_A1_O0),
	.FAB2RAM_A1_O1(Tile_X15Y12_FAB2RAM_A1_O1),
	.FAB2RAM_A1_O2(Tile_X15Y12_FAB2RAM_A1_O2),
	.FAB2RAM_A1_O3(Tile_X15Y12_FAB2RAM_A1_O3),
	.FAB2RAM_C_O0(Tile_X15Y12_FAB2RAM_C_O0),
	.FAB2RAM_C_O1(Tile_X15Y12_FAB2RAM_C_O1),
	.FAB2RAM_C_O2(Tile_X15Y12_FAB2RAM_C_O2),
	.FAB2RAM_C_O3(Tile_X15Y12_FAB2RAM_C_O3),
	.Config_accessC_bit0(Tile_X15Y12_Config_accessC_bit0),
	.Config_accessC_bit1(Tile_X15Y12_Config_accessC_bit1),
	.Config_accessC_bit2(Tile_X15Y12_Config_accessC_bit2),
	.Config_accessC_bit3(Tile_X15Y12_Config_accessC_bit3),
	.UserCLKo(Tile_X15Y12_UserCLKo),
	.FrameData(Tile_X14Y12_FrameData_O), 
	.FrameData_O(Tile_X15Y12_FrameData_O), 
	.FrameStrobe(Tile_X15Y13_FrameStrobe_O),
	.FrameStrobe_O(Tile_X15Y12_FrameStrobe_O)
	);

	S_term_single Tile_X1Y13_S_term_single (
	.S1END(Tile_X1Y12_S1BEG[3:0]),
	.S2MID(Tile_X1Y12_S2BEG[7:0]),
	.S2END(Tile_X1Y12_S2BEGb[7:0]),
	.S4END(Tile_X1Y12_S4BEG[15:0]),
	.SS4END(Tile_X1Y12_SS4BEG[15:0]),
	.N1BEG(Tile_X1Y13_N1BEG[3:0]),
	.N2BEG(Tile_X1Y13_N2BEG[7:0]),
	.N2BEGb(Tile_X1Y13_N2BEGb[7:0]),
	.N4BEG(Tile_X1Y13_N4BEG[15:0]),
	.NN4BEG(Tile_X1Y13_NN4BEG[15:0]),
	.Co(Tile_X1Y13_Co[0:0]),
	.UserCLK(UserCLK),
	.UserCLKo(Tile_X1Y13_UserCLKo),
	.FrameStrobe(Tile_X1_FrameStrobe),
	.FrameStrobe_O(Tile_X1Y13_FrameStrobe_O)
	);

	S_term_single2 Tile_X2Y13_S_term_single2 (
	.S1END(Tile_X2Y12_S1BEG[3:0]),
	.S2MID(Tile_X2Y12_S2BEG[7:0]),
	.S2END(Tile_X2Y12_S2BEGb[7:0]),
	.S4END(Tile_X2Y12_S4BEG[15:0]),
	.SS4END(Tile_X2Y12_SS4BEG[15:0]),
	.N1BEG(Tile_X2Y13_N1BEG[3:0]),
	.N2BEG(Tile_X2Y13_N2BEG[7:0]),
	.N2BEGb(Tile_X2Y13_N2BEGb[7:0]),
	.N4BEG(Tile_X2Y13_N4BEG[15:0]),
	.NN4BEG(Tile_X2Y13_NN4BEG[15:0]),
	.UserCLK(UserCLK),
	.UserCLKo(Tile_X2Y13_UserCLKo),
	.FrameStrobe(Tile_X2_FrameStrobe),
	.FrameStrobe_O(Tile_X2Y13_FrameStrobe_O)
	);

	S_term_single Tile_X3Y13_S_term_single (
	.S1END(Tile_X3Y12_S1BEG[3:0]),
	.S2MID(Tile_X3Y12_S2BEG[7:0]),
	.S2END(Tile_X3Y12_S2BEGb[7:0]),
	.S4END(Tile_X3Y12_S4BEG[15:0]),
	.SS4END(Tile_X3Y12_SS4BEG[15:0]),
	.N1BEG(Tile_X3Y13_N1BEG[3:0]),
	.N2BEG(Tile_X3Y13_N2BEG[7:0]),
	.N2BEGb(Tile_X3Y13_N2BEGb[7:0]),
	.N4BEG(Tile_X3Y13_N4BEG[15:0]),
	.NN4BEG(Tile_X3Y13_NN4BEG[15:0]),
	.Co(Tile_X3Y13_Co[0:0]),
	.UserCLK(UserCLK),
	.UserCLKo(Tile_X3Y13_UserCLKo),
	.FrameStrobe(Tile_X3_FrameStrobe),
	.FrameStrobe_O(Tile_X3Y13_FrameStrobe_O)
	);

	S_term_single Tile_X4Y13_S_term_single (
	.S1END(Tile_X4Y12_S1BEG[3:0]),
	.S2MID(Tile_X4Y12_S2BEG[7:0]),
	.S2END(Tile_X4Y12_S2BEGb[7:0]),
	.S4END(Tile_X4Y12_S4BEG[15:0]),
	.SS4END(Tile_X4Y12_SS4BEG[15:0]),
	.N1BEG(Tile_X4Y13_N1BEG[3:0]),
	.N2BEG(Tile_X4Y13_N2BEG[7:0]),
	.N2BEGb(Tile_X4Y13_N2BEGb[7:0]),
	.N4BEG(Tile_X4Y13_N4BEG[15:0]),
	.NN4BEG(Tile_X4Y13_NN4BEG[15:0]),
	.Co(Tile_X4Y13_Co[0:0]),
	.UserCLK(UserCLK),
	.UserCLKo(Tile_X4Y13_UserCLKo),
	.FrameStrobe(Tile_X4_FrameStrobe),
	.FrameStrobe_O(Tile_X4Y13_FrameStrobe_O)
	);

	S_term_DSP Tile_X5Y13_S_term_DSP (
	.S1END(Tile_X5Y12_S1BEG[3:0]),
	.S2MID(Tile_X5Y12_S2BEG[7:0]),
	.S2END(Tile_X5Y12_S2BEGb[7:0]),
	.S4END(Tile_X5Y12_S4BEG[15:0]),
	.SS4END(Tile_X5Y12_SS4BEG[15:0]),
	.N1BEG(Tile_X5Y13_N1BEG[3:0]),
	.N2BEG(Tile_X5Y13_N2BEG[7:0]),
	.N2BEGb(Tile_X5Y13_N2BEGb[7:0]),
	.N4BEG(Tile_X5Y13_N4BEG[15:0]),
	.NN4BEG(Tile_X5Y13_NN4BEG[15:0]),
	.UserCLK(UserCLK),
	.UserCLKo(Tile_X5Y13_UserCLKo),
	.FrameStrobe(Tile_X5_FrameStrobe),
	.FrameStrobe_O(Tile_X5Y13_FrameStrobe_O)
	);

	S_term_single Tile_X6Y13_S_term_single (
	.S1END(Tile_X6Y12_S1BEG[3:0]),
	.S2MID(Tile_X6Y12_S2BEG[7:0]),
	.S2END(Tile_X6Y12_S2BEGb[7:0]),
	.S4END(Tile_X6Y12_S4BEG[15:0]),
	.SS4END(Tile_X6Y12_SS4BEG[15:0]),
	.N1BEG(Tile_X6Y13_N1BEG[3:0]),
	.N2BEG(Tile_X6Y13_N2BEG[7:0]),
	.N2BEGb(Tile_X6Y13_N2BEGb[7:0]),
	.N4BEG(Tile_X6Y13_N4BEG[15:0]),
	.NN4BEG(Tile_X6Y13_NN4BEG[15:0]),
	.Co(Tile_X6Y13_Co[0:0]),
	.UserCLK(UserCLK),
	.UserCLKo(Tile_X6Y13_UserCLKo),
	.FrameStrobe(Tile_X6_FrameStrobe),
	.FrameStrobe_O(Tile_X6Y13_FrameStrobe_O)
	);

	S_term_single Tile_X7Y13_S_term_single (
	.S1END(Tile_X7Y12_S1BEG[3:0]),
	.S2MID(Tile_X7Y12_S2BEG[7:0]),
	.S2END(Tile_X7Y12_S2BEGb[7:0]),
	.S4END(Tile_X7Y12_S4BEG[15:0]),
	.SS4END(Tile_X7Y12_SS4BEG[15:0]),
	.N1BEG(Tile_X7Y13_N1BEG[3:0]),
	.N2BEG(Tile_X7Y13_N2BEG[7:0]),
	.N2BEGb(Tile_X7Y13_N2BEGb[7:0]),
	.N4BEG(Tile_X7Y13_N4BEG[15:0]),
	.NN4BEG(Tile_X7Y13_NN4BEG[15:0]),
	.Co(Tile_X7Y13_Co[0:0]),
	.UserCLK(UserCLK),
	.UserCLKo(Tile_X7Y13_UserCLKo),
	.FrameStrobe(Tile_X7_FrameStrobe),
	.FrameStrobe_O(Tile_X7Y13_FrameStrobe_O)
	);

	S_term_single Tile_X8Y13_S_term_single (
	.S1END(Tile_X8Y12_S1BEG[3:0]),
	.S2MID(Tile_X8Y12_S2BEG[7:0]),
	.S2END(Tile_X8Y12_S2BEGb[7:0]),
	.S4END(Tile_X8Y12_S4BEG[15:0]),
	.SS4END(Tile_X8Y12_SS4BEG[15:0]),
	.N1BEG(Tile_X8Y13_N1BEG[3:0]),
	.N2BEG(Tile_X8Y13_N2BEG[7:0]),
	.N2BEGb(Tile_X8Y13_N2BEGb[7:0]),
	.N4BEG(Tile_X8Y13_N4BEG[15:0]),
	.NN4BEG(Tile_X8Y13_NN4BEG[15:0]),
	.Co(Tile_X8Y13_Co[0:0]),
	.UserCLK(UserCLK),
	.UserCLKo(Tile_X8Y13_UserCLKo),
	.FrameStrobe(Tile_X8_FrameStrobe),
	.FrameStrobe_O(Tile_X8Y13_FrameStrobe_O)
	);

	S_term_DSP Tile_X9Y13_S_term_DSP (
	.S1END(Tile_X9Y12_S1BEG[3:0]),
	.S2MID(Tile_X9Y12_S2BEG[7:0]),
	.S2END(Tile_X9Y12_S2BEGb[7:0]),
	.S4END(Tile_X9Y12_S4BEG[15:0]),
	.SS4END(Tile_X9Y12_SS4BEG[15:0]),
	.N1BEG(Tile_X9Y13_N1BEG[3:0]),
	.N2BEG(Tile_X9Y13_N2BEG[7:0]),
	.N2BEGb(Tile_X9Y13_N2BEGb[7:0]),
	.N4BEG(Tile_X9Y13_N4BEG[15:0]),
	.NN4BEG(Tile_X9Y13_NN4BEG[15:0]),
	.UserCLK(UserCLK),
	.UserCLKo(Tile_X9Y13_UserCLKo),
	.FrameStrobe(Tile_X9_FrameStrobe),
	.FrameStrobe_O(Tile_X9Y13_FrameStrobe_O)
	);

	S_term_single Tile_X10Y13_S_term_single (
	.S1END(Tile_X10Y12_S1BEG[3:0]),
	.S2MID(Tile_X10Y12_S2BEG[7:0]),
	.S2END(Tile_X10Y12_S2BEGb[7:0]),
	.S4END(Tile_X10Y12_S4BEG[15:0]),
	.SS4END(Tile_X10Y12_SS4BEG[15:0]),
	.N1BEG(Tile_X10Y13_N1BEG[3:0]),
	.N2BEG(Tile_X10Y13_N2BEG[7:0]),
	.N2BEGb(Tile_X10Y13_N2BEGb[7:0]),
	.N4BEG(Tile_X10Y13_N4BEG[15:0]),
	.NN4BEG(Tile_X10Y13_NN4BEG[15:0]),
	.Co(Tile_X10Y13_Co[0:0]),
	.UserCLK(UserCLK),
	.UserCLKo(Tile_X10Y13_UserCLKo),
	.FrameStrobe(Tile_X10_FrameStrobe),
	.FrameStrobe_O(Tile_X10Y13_FrameStrobe_O)
	);

	S_term_single Tile_X11Y13_S_term_single (
	.S1END(Tile_X11Y12_S1BEG[3:0]),
	.S2MID(Tile_X11Y12_S2BEG[7:0]),
	.S2END(Tile_X11Y12_S2BEGb[7:0]),
	.S4END(Tile_X11Y12_S4BEG[15:0]),
	.SS4END(Tile_X11Y12_SS4BEG[15:0]),
	.N1BEG(Tile_X11Y13_N1BEG[3:0]),
	.N2BEG(Tile_X11Y13_N2BEG[7:0]),
	.N2BEGb(Tile_X11Y13_N2BEGb[7:0]),
	.N4BEG(Tile_X11Y13_N4BEG[15:0]),
	.NN4BEG(Tile_X11Y13_NN4BEG[15:0]),
	.Co(Tile_X11Y13_Co[0:0]),
	.UserCLK(UserCLK),
	.UserCLKo(Tile_X11Y13_UserCLKo),
	.FrameStrobe(Tile_X11_FrameStrobe),
	.FrameStrobe_O(Tile_X11Y13_FrameStrobe_O)
	);

	S_term_single Tile_X12Y13_S_term_single (
	.S1END(Tile_X12Y12_S1BEG[3:0]),
	.S2MID(Tile_X12Y12_S2BEG[7:0]),
	.S2END(Tile_X12Y12_S2BEGb[7:0]),
	.S4END(Tile_X12Y12_S4BEG[15:0]),
	.SS4END(Tile_X12Y12_SS4BEG[15:0]),
	.N1BEG(Tile_X12Y13_N1BEG[3:0]),
	.N2BEG(Tile_X12Y13_N2BEG[7:0]),
	.N2BEGb(Tile_X12Y13_N2BEGb[7:0]),
	.N4BEG(Tile_X12Y13_N4BEG[15:0]),
	.NN4BEG(Tile_X12Y13_NN4BEG[15:0]),
	.Co(Tile_X12Y13_Co[0:0]),
	.UserCLK(UserCLK),
	.UserCLKo(Tile_X12Y13_UserCLKo),
	.FrameStrobe(Tile_X12_FrameStrobe),
	.FrameStrobe_O(Tile_X12Y13_FrameStrobe_O)
	);

	S_term_single2 Tile_X13Y13_S_term_single2 (
	.S1END(Tile_X13Y12_S1BEG[3:0]),
	.S2MID(Tile_X13Y12_S2BEG[7:0]),
	.S2END(Tile_X13Y12_S2BEGb[7:0]),
	.S4END(Tile_X13Y12_S4BEG[15:0]),
	.SS4END(Tile_X13Y12_SS4BEG[15:0]),
	.N1BEG(Tile_X13Y13_N1BEG[3:0]),
	.N2BEG(Tile_X13Y13_N2BEG[7:0]),
	.N2BEGb(Tile_X13Y13_N2BEGb[7:0]),
	.N4BEG(Tile_X13Y13_N4BEG[15:0]),
	.NN4BEG(Tile_X13Y13_NN4BEG[15:0]),
	.UserCLK(UserCLK),
	.UserCLKo(Tile_X13Y13_UserCLKo),
	.FrameStrobe(Tile_X13_FrameStrobe),
	.FrameStrobe_O(Tile_X13Y13_FrameStrobe_O)
	);

	S_term_single Tile_X14Y13_S_term_single (
	.S1END(Tile_X14Y12_S1BEG[3:0]),
	.S2MID(Tile_X14Y12_S2BEG[7:0]),
	.S2END(Tile_X14Y12_S2BEGb[7:0]),
	.S4END(Tile_X14Y12_S4BEG[15:0]),
	.SS4END(Tile_X14Y12_SS4BEG[15:0]),
	.N1BEG(Tile_X14Y13_N1BEG[3:0]),
	.N2BEG(Tile_X14Y13_N2BEG[7:0]),
	.N2BEGb(Tile_X14Y13_N2BEGb[7:0]),
	.N4BEG(Tile_X14Y13_N4BEG[15:0]),
	.NN4BEG(Tile_X14Y13_NN4BEG[15:0]),
	.Co(Tile_X14Y13_Co[0:0]),
	.UserCLK(UserCLK),
	.UserCLKo(Tile_X14Y13_UserCLKo),
	.FrameStrobe(Tile_X14_FrameStrobe),
	.FrameStrobe_O(Tile_X14Y13_FrameStrobe_O)
	);

	S_term_RAM_IO Tile_X15Y13_S_term_RAM_IO (
	.S1END(Tile_X15Y12_S1BEG[3:0]),
	.S2MID(Tile_X15Y12_S2BEG[7:0]),
	.S2END(Tile_X15Y12_S2BEGb[7:0]),
	.S4END(Tile_X15Y12_S4BEG[15:0]),
	.N1BEG(Tile_X15Y13_N1BEG[3:0]),
	.N2BEG(Tile_X15Y13_N2BEG[7:0]),
	.N2BEGb(Tile_X15Y13_N2BEGb[7:0]),
	.N4BEG(Tile_X15Y13_N4BEG[15:0]),
	.UserCLK(UserCLK),
	.UserCLKo(Tile_X15Y13_UserCLKo),
	.FrameStrobe(Tile_X15_FrameStrobe),
	.FrameStrobe_O(Tile_X15Y13_FrameStrobe_O)
	);


	DSP Tile_X5Y1_X5Y2_DSP_tile (
	.top_E1END(Tile_X4Y1_E1BEG[3:0]),
	.top_E2MID(Tile_X4Y1_E2BEG[7:0]),
	.top_E2END(Tile_X4Y1_E2BEGb[7:0]),
	.top_EE4END(Tile_X4Y1_EE4BEG[15:0]),
	.top_E6END(Tile_X4Y1_E6BEG[11:0]),
	.top_S1END(Tile_X5Y0_S1BEG[3:0]),
	.top_S2MID(Tile_X5Y0_S2BEG[7:0]),
	.top_S2END(Tile_X5Y0_S2BEGb[7:0]),
	.top_S4END(Tile_X5Y0_S4BEG[15:0]),
	.top_SS4END(Tile_X5Y0_SS4BEG[15:0]),
	.top_W1END(Tile_X6Y1_W1BEG[3:0]),
	.top_W2MID(Tile_X6Y1_W2BEG[7:0]),
	.top_W2END(Tile_X6Y1_W2BEGb[7:0]),
	.top_WW4END(Tile_X6Y1_WW4BEG[15:0]),
	.top_W6END(Tile_X6Y1_W6BEG[11:0]),
	.top_N1BEG(Tile_X5Y1_N1BEG[3:0]),
	.top_N2BEG(Tile_X5Y1_N2BEG[7:0]),
	.top_N2BEGb(Tile_X5Y1_N2BEGb[7:0]),
	.top_N4BEG(Tile_X5Y1_N4BEG[15:0]),
	.top_NN4BEG(Tile_X5Y1_NN4BEG[15:0]),
	.top_E1BEG(Tile_X5Y1_E1BEG[3:0]),
	.top_E2BEG(Tile_X5Y1_E2BEG[7:0]),
	.top_E2BEGb(Tile_X5Y1_E2BEGb[7:0]),
	.top_EE4BEG(Tile_X5Y1_EE4BEG[15:0]),
	.top_E6BEG(Tile_X5Y1_E6BEG[11:0]),
	.top_W1BEG(Tile_X5Y1_W1BEG[3:0]),
	.top_W2BEG(Tile_X5Y1_W2BEG[7:0]),
	.top_W2BEGb(Tile_X5Y1_W2BEGb[7:0]),
	.top_WW4BEG(Tile_X5Y1_WW4BEG[15:0]),
	.top_W6BEG(Tile_X5Y1_W6BEG[11:0]),
	.top_FrameData(Tile_X4Y1_FrameData_O),
	.top_FrameData_O(Tile_X5Y1_FrameData_O),
	.FrameStrobe_O(Tile_X5Y1_FrameStrobe_O),
	.UserCLKo(Tile_X5Y1_UserCLKo),
	.bot_N1END(Tile_X5Y3_N1BEG[3:0]),
	.bot_N2MID(Tile_X5Y3_N2BEG[7:0]),
	.bot_N2END(Tile_X5Y3_N2BEGb[7:0]),
	.bot_N4END(Tile_X5Y3_N4BEG[15:0]),
	.bot_NN4END(Tile_X5Y3_NN4BEG[15:0]),
	.bot_E1END(Tile_X4Y2_E1BEG[3:0]),
	.bot_E2MID(Tile_X4Y2_E2BEG[7:0]),
	.bot_E2END(Tile_X4Y2_E2BEGb[7:0]),
	.bot_EE4END(Tile_X4Y2_EE4BEG[15:0]),
	.bot_E6END(Tile_X4Y2_E6BEG[11:0]),
	.bot_W1END(Tile_X6Y2_W1BEG[3:0]),
	.bot_W2MID(Tile_X6Y2_W2BEG[7:0]),
	.bot_W2END(Tile_X6Y2_W2BEGb[7:0]),
	.bot_WW4END(Tile_X6Y2_WW4BEG[15:0]),
	.bot_W6END(Tile_X6Y2_W6BEG[11:0]),
	.bot_E1BEG(Tile_X5Y2_E1BEG[3:0]),
	.bot_E2BEG(Tile_X5Y2_E2BEG[7:0]),
	.bot_E2BEGb(Tile_X5Y2_E2BEGb[7:0]),
	.bot_EE4BEG(Tile_X5Y2_EE4BEG[15:0]),
	.bot_E6BEG(Tile_X5Y2_E6BEG[11:0]),
	.bot_S1BEG(Tile_X5Y2_S1BEG[3:0]),
	.bot_S2BEG(Tile_X5Y2_S2BEG[7:0]),
	.bot_S2BEGb(Tile_X5Y2_S2BEGb[7:0]),
	.bot_S4BEG(Tile_X5Y2_S4BEG[15:0]),
	.bot_SS4BEG(Tile_X5Y2_SS4BEG[15:0]),
	.bot_W1BEG(Tile_X5Y2_W1BEG[3:0]),
	.bot_W2BEG(Tile_X5Y2_W2BEG[7:0]),
	.bot_W2BEGb(Tile_X5Y2_W2BEGb[7:0]),
	.bot_WW4BEG(Tile_X5Y2_WW4BEG[15:0]),
	.bot_W6BEG(Tile_X5Y2_W6BEG[11:0]),
	.UserCLK(Tile_X5Y3_UserCLKo),
	.bot_FrameData(Tile_X4Y2_FrameData_O),
	.bot_FrameData_O(Tile_X5Y2_FrameData_O),
	.FrameStrobe(Tile_X5Y3_FrameStrobe_O)
	);

	DSP Tile_X9Y1_X9Y2_DSP_tile (
	.top_E1END(Tile_X8Y1_E1BEG[3:0]),
	.top_E2MID(Tile_X8Y1_E2BEG[7:0]),
	.top_E2END(Tile_X8Y1_E2BEGb[7:0]),
	.top_EE4END(Tile_X8Y1_EE4BEG[15:0]),
	.top_E6END(Tile_X8Y1_E6BEG[11:0]),
	.top_S1END(Tile_X9Y0_S1BEG[3:0]),
	.top_S2MID(Tile_X9Y0_S2BEG[7:0]),
	.top_S2END(Tile_X9Y0_S2BEGb[7:0]),
	.top_S4END(Tile_X9Y0_S4BEG[15:0]),
	.top_SS4END(Tile_X9Y0_SS4BEG[15:0]),
	.top_W1END(Tile_X10Y1_W1BEG[3:0]),
	.top_W2MID(Tile_X10Y1_W2BEG[7:0]),
	.top_W2END(Tile_X10Y1_W2BEGb[7:0]),
	.top_WW4END(Tile_X10Y1_WW4BEG[15:0]),
	.top_W6END(Tile_X10Y1_W6BEG[11:0]),
	.top_N1BEG(Tile_X9Y1_N1BEG[3:0]),
	.top_N2BEG(Tile_X9Y1_N2BEG[7:0]),
	.top_N2BEGb(Tile_X9Y1_N2BEGb[7:0]),
	.top_N4BEG(Tile_X9Y1_N4BEG[15:0]),
	.top_NN4BEG(Tile_X9Y1_NN4BEG[15:0]),
	.top_E1BEG(Tile_X9Y1_E1BEG[3:0]),
	.top_E2BEG(Tile_X9Y1_E2BEG[7:0]),
	.top_E2BEGb(Tile_X9Y1_E2BEGb[7:0]),
	.top_EE4BEG(Tile_X9Y1_EE4BEG[15:0]),
	.top_E6BEG(Tile_X9Y1_E6BEG[11:0]),
	.top_W1BEG(Tile_X9Y1_W1BEG[3:0]),
	.top_W2BEG(Tile_X9Y1_W2BEG[7:0]),
	.top_W2BEGb(Tile_X9Y1_W2BEGb[7:0]),
	.top_WW4BEG(Tile_X9Y1_WW4BEG[15:0]),
	.top_W6BEG(Tile_X9Y1_W6BEG[11:0]),
	.top_FrameData(Tile_X8Y1_FrameData_O),
	.top_FrameData_O(Tile_X9Y1_FrameData_O),
	.FrameStrobe_O(Tile_X9Y1_FrameStrobe_O),
	.UserCLKo(Tile_X9Y1_UserCLKo),
	.bot_N1END(Tile_X9Y3_N1BEG[3:0]),
	.bot_N2MID(Tile_X9Y3_N2BEG[7:0]),
	.bot_N2END(Tile_X9Y3_N2BEGb[7:0]),
	.bot_N4END(Tile_X9Y3_N4BEG[15:0]),
	.bot_NN4END(Tile_X9Y3_NN4BEG[15:0]),
	.bot_E1END(Tile_X8Y2_E1BEG[3:0]),
	.bot_E2MID(Tile_X8Y2_E2BEG[7:0]),
	.bot_E2END(Tile_X8Y2_E2BEGb[7:0]),
	.bot_EE4END(Tile_X8Y2_EE4BEG[15:0]),
	.bot_E6END(Tile_X8Y2_E6BEG[11:0]),
	.bot_W1END(Tile_X10Y2_W1BEG[3:0]),
	.bot_W2MID(Tile_X10Y2_W2BEG[7:0]),
	.bot_W2END(Tile_X10Y2_W2BEGb[7:0]),
	.bot_WW4END(Tile_X10Y2_WW4BEG[15:0]),
	.bot_W6END(Tile_X10Y2_W6BEG[11:0]),
	.bot_E1BEG(Tile_X9Y2_E1BEG[3:0]),
	.bot_E2BEG(Tile_X9Y2_E2BEG[7:0]),
	.bot_E2BEGb(Tile_X9Y2_E2BEGb[7:0]),
	.bot_EE4BEG(Tile_X9Y2_EE4BEG[15:0]),
	.bot_E6BEG(Tile_X9Y2_E6BEG[11:0]),
	.bot_S1BEG(Tile_X9Y2_S1BEG[3:0]),
	.bot_S2BEG(Tile_X9Y2_S2BEG[7:0]),
	.bot_S2BEGb(Tile_X9Y2_S2BEGb[7:0]),
	.bot_S4BEG(Tile_X9Y2_S4BEG[15:0]),
	.bot_SS4BEG(Tile_X9Y2_SS4BEG[15:0]),
	.bot_W1BEG(Tile_X9Y2_W1BEG[3:0]),
	.bot_W2BEG(Tile_X9Y2_W2BEG[7:0]),
	.bot_W2BEGb(Tile_X9Y2_W2BEGb[7:0]),
	.bot_WW4BEG(Tile_X9Y2_WW4BEG[15:0]),
	.bot_W6BEG(Tile_X9Y2_W6BEG[11:0]),
	.UserCLK(Tile_X9Y3_UserCLKo),
	.bot_FrameData(Tile_X8Y2_FrameData_O),
	.bot_FrameData_O(Tile_X9Y2_FrameData_O),
	.FrameStrobe(Tile_X9Y3_FrameStrobe_O)
	);

	DSP Tile_X5Y3_X5Y4_DSP_tile (
	.top_E1END(Tile_X4Y3_E1BEG[3:0]),
	.top_E2MID(Tile_X4Y3_E2BEG[7:0]),
	.top_E2END(Tile_X4Y3_E2BEGb[7:0]),
	.top_EE4END(Tile_X4Y3_EE4BEG[15:0]),
	.top_E6END(Tile_X4Y3_E6BEG[11:0]),
	.top_S1END(Tile_X5Y2_S1BEG[3:0]),
	.top_S2MID(Tile_X5Y2_S2BEG[7:0]),
	.top_S2END(Tile_X5Y2_S2BEGb[7:0]),
	.top_S4END(Tile_X5Y2_S4BEG[15:0]),
	.top_SS4END(Tile_X5Y2_SS4BEG[15:0]),
	.top_W1END(Tile_X6Y3_W1BEG[3:0]),
	.top_W2MID(Tile_X6Y3_W2BEG[7:0]),
	.top_W2END(Tile_X6Y3_W2BEGb[7:0]),
	.top_WW4END(Tile_X6Y3_WW4BEG[15:0]),
	.top_W6END(Tile_X6Y3_W6BEG[11:0]),
	.top_N1BEG(Tile_X5Y3_N1BEG[3:0]),
	.top_N2BEG(Tile_X5Y3_N2BEG[7:0]),
	.top_N2BEGb(Tile_X5Y3_N2BEGb[7:0]),
	.top_N4BEG(Tile_X5Y3_N4BEG[15:0]),
	.top_NN4BEG(Tile_X5Y3_NN4BEG[15:0]),
	.top_E1BEG(Tile_X5Y3_E1BEG[3:0]),
	.top_E2BEG(Tile_X5Y3_E2BEG[7:0]),
	.top_E2BEGb(Tile_X5Y3_E2BEGb[7:0]),
	.top_EE4BEG(Tile_X5Y3_EE4BEG[15:0]),
	.top_E6BEG(Tile_X5Y3_E6BEG[11:0]),
	.top_W1BEG(Tile_X5Y3_W1BEG[3:0]),
	.top_W2BEG(Tile_X5Y3_W2BEG[7:0]),
	.top_W2BEGb(Tile_X5Y3_W2BEGb[7:0]),
	.top_WW4BEG(Tile_X5Y3_WW4BEG[15:0]),
	.top_W6BEG(Tile_X5Y3_W6BEG[11:0]),
	.top_FrameData(Tile_X4Y3_FrameData_O),
	.top_FrameData_O(Tile_X5Y3_FrameData_O),
	.FrameStrobe_O(Tile_X5Y3_FrameStrobe_O),
	.UserCLKo(Tile_X5Y3_UserCLKo),
	.bot_N1END(Tile_X5Y5_N1BEG[3:0]),
	.bot_N2MID(Tile_X5Y5_N2BEG[7:0]),
	.bot_N2END(Tile_X5Y5_N2BEGb[7:0]),
	.bot_N4END(Tile_X5Y5_N4BEG[15:0]),
	.bot_NN4END(Tile_X5Y5_NN4BEG[15:0]),
	.bot_E1END(Tile_X4Y4_E1BEG[3:0]),
	.bot_E2MID(Tile_X4Y4_E2BEG[7:0]),
	.bot_E2END(Tile_X4Y4_E2BEGb[7:0]),
	.bot_EE4END(Tile_X4Y4_EE4BEG[15:0]),
	.bot_E6END(Tile_X4Y4_E6BEG[11:0]),
	.bot_W1END(Tile_X6Y4_W1BEG[3:0]),
	.bot_W2MID(Tile_X6Y4_W2BEG[7:0]),
	.bot_W2END(Tile_X6Y4_W2BEGb[7:0]),
	.bot_WW4END(Tile_X6Y4_WW4BEG[15:0]),
	.bot_W6END(Tile_X6Y4_W6BEG[11:0]),
	.bot_E1BEG(Tile_X5Y4_E1BEG[3:0]),
	.bot_E2BEG(Tile_X5Y4_E2BEG[7:0]),
	.bot_E2BEGb(Tile_X5Y4_E2BEGb[7:0]),
	.bot_EE4BEG(Tile_X5Y4_EE4BEG[15:0]),
	.bot_E6BEG(Tile_X5Y4_E6BEG[11:0]),
	.bot_S1BEG(Tile_X5Y4_S1BEG[3:0]),
	.bot_S2BEG(Tile_X5Y4_S2BEG[7:0]),
	.bot_S2BEGb(Tile_X5Y4_S2BEGb[7:0]),
	.bot_S4BEG(Tile_X5Y4_S4BEG[15:0]),
	.bot_SS4BEG(Tile_X5Y4_SS4BEG[15:0]),
	.bot_W1BEG(Tile_X5Y4_W1BEG[3:0]),
	.bot_W2BEG(Tile_X5Y4_W2BEG[7:0]),
	.bot_W2BEGb(Tile_X5Y4_W2BEGb[7:0]),
	.bot_WW4BEG(Tile_X5Y4_WW4BEG[15:0]),
	.bot_W6BEG(Tile_X5Y4_W6BEG[11:0]),
	.UserCLK(Tile_X5Y5_UserCLKo),
	.bot_FrameData(Tile_X4Y4_FrameData_O),
	.bot_FrameData_O(Tile_X5Y4_FrameData_O),
	.FrameStrobe(Tile_X5Y5_FrameStrobe_O)
	);

	DSP Tile_X9Y3_X9Y4_DSP_tile (
	.top_E1END(Tile_X8Y3_E1BEG[3:0]),
	.top_E2MID(Tile_X8Y3_E2BEG[7:0]),
	.top_E2END(Tile_X8Y3_E2BEGb[7:0]),
	.top_EE4END(Tile_X8Y3_EE4BEG[15:0]),
	.top_E6END(Tile_X8Y3_E6BEG[11:0]),
	.top_S1END(Tile_X9Y2_S1BEG[3:0]),
	.top_S2MID(Tile_X9Y2_S2BEG[7:0]),
	.top_S2END(Tile_X9Y2_S2BEGb[7:0]),
	.top_S4END(Tile_X9Y2_S4BEG[15:0]),
	.top_SS4END(Tile_X9Y2_SS4BEG[15:0]),
	.top_W1END(Tile_X10Y3_W1BEG[3:0]),
	.top_W2MID(Tile_X10Y3_W2BEG[7:0]),
	.top_W2END(Tile_X10Y3_W2BEGb[7:0]),
	.top_WW4END(Tile_X10Y3_WW4BEG[15:0]),
	.top_W6END(Tile_X10Y3_W6BEG[11:0]),
	.top_N1BEG(Tile_X9Y3_N1BEG[3:0]),
	.top_N2BEG(Tile_X9Y3_N2BEG[7:0]),
	.top_N2BEGb(Tile_X9Y3_N2BEGb[7:0]),
	.top_N4BEG(Tile_X9Y3_N4BEG[15:0]),
	.top_NN4BEG(Tile_X9Y3_NN4BEG[15:0]),
	.top_E1BEG(Tile_X9Y3_E1BEG[3:0]),
	.top_E2BEG(Tile_X9Y3_E2BEG[7:0]),
	.top_E2BEGb(Tile_X9Y3_E2BEGb[7:0]),
	.top_EE4BEG(Tile_X9Y3_EE4BEG[15:0]),
	.top_E6BEG(Tile_X9Y3_E6BEG[11:0]),
	.top_W1BEG(Tile_X9Y3_W1BEG[3:0]),
	.top_W2BEG(Tile_X9Y3_W2BEG[7:0]),
	.top_W2BEGb(Tile_X9Y3_W2BEGb[7:0]),
	.top_WW4BEG(Tile_X9Y3_WW4BEG[15:0]),
	.top_W6BEG(Tile_X9Y3_W6BEG[11:0]),
	.top_FrameData(Tile_X8Y3_FrameData_O),
	.top_FrameData_O(Tile_X9Y3_FrameData_O),
	.FrameStrobe_O(Tile_X9Y3_FrameStrobe_O),
	.UserCLKo(Tile_X9Y3_UserCLKo),
	.bot_N1END(Tile_X9Y5_N1BEG[3:0]),
	.bot_N2MID(Tile_X9Y5_N2BEG[7:0]),
	.bot_N2END(Tile_X9Y5_N2BEGb[7:0]),
	.bot_N4END(Tile_X9Y5_N4BEG[15:0]),
	.bot_NN4END(Tile_X9Y5_NN4BEG[15:0]),
	.bot_E1END(Tile_X8Y4_E1BEG[3:0]),
	.bot_E2MID(Tile_X8Y4_E2BEG[7:0]),
	.bot_E2END(Tile_X8Y4_E2BEGb[7:0]),
	.bot_EE4END(Tile_X8Y4_EE4BEG[15:0]),
	.bot_E6END(Tile_X8Y4_E6BEG[11:0]),
	.bot_W1END(Tile_X10Y4_W1BEG[3:0]),
	.bot_W2MID(Tile_X10Y4_W2BEG[7:0]),
	.bot_W2END(Tile_X10Y4_W2BEGb[7:0]),
	.bot_WW4END(Tile_X10Y4_WW4BEG[15:0]),
	.bot_W6END(Tile_X10Y4_W6BEG[11:0]),
	.bot_E1BEG(Tile_X9Y4_E1BEG[3:0]),
	.bot_E2BEG(Tile_X9Y4_E2BEG[7:0]),
	.bot_E2BEGb(Tile_X9Y4_E2BEGb[7:0]),
	.bot_EE4BEG(Tile_X9Y4_EE4BEG[15:0]),
	.bot_E6BEG(Tile_X9Y4_E6BEG[11:0]),
	.bot_S1BEG(Tile_X9Y4_S1BEG[3:0]),
	.bot_S2BEG(Tile_X9Y4_S2BEG[7:0]),
	.bot_S2BEGb(Tile_X9Y4_S2BEGb[7:0]),
	.bot_S4BEG(Tile_X9Y4_S4BEG[15:0]),
	.bot_SS4BEG(Tile_X9Y4_SS4BEG[15:0]),
	.bot_W1BEG(Tile_X9Y4_W1BEG[3:0]),
	.bot_W2BEG(Tile_X9Y4_W2BEG[7:0]),
	.bot_W2BEGb(Tile_X9Y4_W2BEGb[7:0]),
	.bot_WW4BEG(Tile_X9Y4_WW4BEG[15:0]),
	.bot_W6BEG(Tile_X9Y4_W6BEG[11:0]),
	.UserCLK(Tile_X9Y5_UserCLKo),
	.bot_FrameData(Tile_X8Y4_FrameData_O),
	.bot_FrameData_O(Tile_X9Y4_FrameData_O),
	.FrameStrobe(Tile_X9Y5_FrameStrobe_O)
	);

	DSP Tile_X5Y5_X5Y6_DSP_tile (
	.top_E1END(Tile_X4Y5_E1BEG[3:0]),
	.top_E2MID(Tile_X4Y5_E2BEG[7:0]),
	.top_E2END(Tile_X4Y5_E2BEGb[7:0]),
	.top_EE4END(Tile_X4Y5_EE4BEG[15:0]),
	.top_E6END(Tile_X4Y5_E6BEG[11:0]),
	.top_S1END(Tile_X5Y4_S1BEG[3:0]),
	.top_S2MID(Tile_X5Y4_S2BEG[7:0]),
	.top_S2END(Tile_X5Y4_S2BEGb[7:0]),
	.top_S4END(Tile_X5Y4_S4BEG[15:0]),
	.top_SS4END(Tile_X5Y4_SS4BEG[15:0]),
	.top_W1END(Tile_X6Y5_W1BEG[3:0]),
	.top_W2MID(Tile_X6Y5_W2BEG[7:0]),
	.top_W2END(Tile_X6Y5_W2BEGb[7:0]),
	.top_WW4END(Tile_X6Y5_WW4BEG[15:0]),
	.top_W6END(Tile_X6Y5_W6BEG[11:0]),
	.top_N1BEG(Tile_X5Y5_N1BEG[3:0]),
	.top_N2BEG(Tile_X5Y5_N2BEG[7:0]),
	.top_N2BEGb(Tile_X5Y5_N2BEGb[7:0]),
	.top_N4BEG(Tile_X5Y5_N4BEG[15:0]),
	.top_NN4BEG(Tile_X5Y5_NN4BEG[15:0]),
	.top_E1BEG(Tile_X5Y5_E1BEG[3:0]),
	.top_E2BEG(Tile_X5Y5_E2BEG[7:0]),
	.top_E2BEGb(Tile_X5Y5_E2BEGb[7:0]),
	.top_EE4BEG(Tile_X5Y5_EE4BEG[15:0]),
	.top_E6BEG(Tile_X5Y5_E6BEG[11:0]),
	.top_W1BEG(Tile_X5Y5_W1BEG[3:0]),
	.top_W2BEG(Tile_X5Y5_W2BEG[7:0]),
	.top_W2BEGb(Tile_X5Y5_W2BEGb[7:0]),
	.top_WW4BEG(Tile_X5Y5_WW4BEG[15:0]),
	.top_W6BEG(Tile_X5Y5_W6BEG[11:0]),
	.top_FrameData(Tile_X4Y5_FrameData_O),
	.top_FrameData_O(Tile_X5Y5_FrameData_O),
	.FrameStrobe_O(Tile_X5Y5_FrameStrobe_O),
	.UserCLKo(Tile_X5Y5_UserCLKo),
	.bot_N1END(Tile_X5Y7_N1BEG[3:0]),
	.bot_N2MID(Tile_X5Y7_N2BEG[7:0]),
	.bot_N2END(Tile_X5Y7_N2BEGb[7:0]),
	.bot_N4END(Tile_X5Y7_N4BEG[15:0]),
	.bot_NN4END(Tile_X5Y7_NN4BEG[15:0]),
	.bot_E1END(Tile_X4Y6_E1BEG[3:0]),
	.bot_E2MID(Tile_X4Y6_E2BEG[7:0]),
	.bot_E2END(Tile_X4Y6_E2BEGb[7:0]),
	.bot_EE4END(Tile_X4Y6_EE4BEG[15:0]),
	.bot_E6END(Tile_X4Y6_E6BEG[11:0]),
	.bot_W1END(Tile_X6Y6_W1BEG[3:0]),
	.bot_W2MID(Tile_X6Y6_W2BEG[7:0]),
	.bot_W2END(Tile_X6Y6_W2BEGb[7:0]),
	.bot_WW4END(Tile_X6Y6_WW4BEG[15:0]),
	.bot_W6END(Tile_X6Y6_W6BEG[11:0]),
	.bot_E1BEG(Tile_X5Y6_E1BEG[3:0]),
	.bot_E2BEG(Tile_X5Y6_E2BEG[7:0]),
	.bot_E2BEGb(Tile_X5Y6_E2BEGb[7:0]),
	.bot_EE4BEG(Tile_X5Y6_EE4BEG[15:0]),
	.bot_E6BEG(Tile_X5Y6_E6BEG[11:0]),
	.bot_S1BEG(Tile_X5Y6_S1BEG[3:0]),
	.bot_S2BEG(Tile_X5Y6_S2BEG[7:0]),
	.bot_S2BEGb(Tile_X5Y6_S2BEGb[7:0]),
	.bot_S4BEG(Tile_X5Y6_S4BEG[15:0]),
	.bot_SS4BEG(Tile_X5Y6_SS4BEG[15:0]),
	.bot_W1BEG(Tile_X5Y6_W1BEG[3:0]),
	.bot_W2BEG(Tile_X5Y6_W2BEG[7:0]),
	.bot_W2BEGb(Tile_X5Y6_W2BEGb[7:0]),
	.bot_WW4BEG(Tile_X5Y6_WW4BEG[15:0]),
	.bot_W6BEG(Tile_X5Y6_W6BEG[11:0]),
	.UserCLK(Tile_X5Y7_UserCLKo),
	.bot_FrameData(Tile_X4Y6_FrameData_O),
	.bot_FrameData_O(Tile_X5Y6_FrameData_O),
	.FrameStrobe(Tile_X5Y7_FrameStrobe_O)
	);

	DSP Tile_X9Y5_X9Y6_DSP_tile (
	.top_E1END(Tile_X8Y5_E1BEG[3:0]),
	.top_E2MID(Tile_X8Y5_E2BEG[7:0]),
	.top_E2END(Tile_X8Y5_E2BEGb[7:0]),
	.top_EE4END(Tile_X8Y5_EE4BEG[15:0]),
	.top_E6END(Tile_X8Y5_E6BEG[11:0]),
	.top_S1END(Tile_X9Y4_S1BEG[3:0]),
	.top_S2MID(Tile_X9Y4_S2BEG[7:0]),
	.top_S2END(Tile_X9Y4_S2BEGb[7:0]),
	.top_S4END(Tile_X9Y4_S4BEG[15:0]),
	.top_SS4END(Tile_X9Y4_SS4BEG[15:0]),
	.top_W1END(Tile_X10Y5_W1BEG[3:0]),
	.top_W2MID(Tile_X10Y5_W2BEG[7:0]),
	.top_W2END(Tile_X10Y5_W2BEGb[7:0]),
	.top_WW4END(Tile_X10Y5_WW4BEG[15:0]),
	.top_W6END(Tile_X10Y5_W6BEG[11:0]),
	.top_N1BEG(Tile_X9Y5_N1BEG[3:0]),
	.top_N2BEG(Tile_X9Y5_N2BEG[7:0]),
	.top_N2BEGb(Tile_X9Y5_N2BEGb[7:0]),
	.top_N4BEG(Tile_X9Y5_N4BEG[15:0]),
	.top_NN4BEG(Tile_X9Y5_NN4BEG[15:0]),
	.top_E1BEG(Tile_X9Y5_E1BEG[3:0]),
	.top_E2BEG(Tile_X9Y5_E2BEG[7:0]),
	.top_E2BEGb(Tile_X9Y5_E2BEGb[7:0]),
	.top_EE4BEG(Tile_X9Y5_EE4BEG[15:0]),
	.top_E6BEG(Tile_X9Y5_E6BEG[11:0]),
	.top_W1BEG(Tile_X9Y5_W1BEG[3:0]),
	.top_W2BEG(Tile_X9Y5_W2BEG[7:0]),
	.top_W2BEGb(Tile_X9Y5_W2BEGb[7:0]),
	.top_WW4BEG(Tile_X9Y5_WW4BEG[15:0]),
	.top_W6BEG(Tile_X9Y5_W6BEG[11:0]),
	.top_FrameData(Tile_X8Y5_FrameData_O),
	.top_FrameData_O(Tile_X9Y5_FrameData_O),
	.FrameStrobe_O(Tile_X9Y5_FrameStrobe_O),
	.UserCLKo(Tile_X9Y5_UserCLKo),
	.bot_N1END(Tile_X9Y7_N1BEG[3:0]),
	.bot_N2MID(Tile_X9Y7_N2BEG[7:0]),
	.bot_N2END(Tile_X9Y7_N2BEGb[7:0]),
	.bot_N4END(Tile_X9Y7_N4BEG[15:0]),
	.bot_NN4END(Tile_X9Y7_NN4BEG[15:0]),
	.bot_E1END(Tile_X8Y6_E1BEG[3:0]),
	.bot_E2MID(Tile_X8Y6_E2BEG[7:0]),
	.bot_E2END(Tile_X8Y6_E2BEGb[7:0]),
	.bot_EE4END(Tile_X8Y6_EE4BEG[15:0]),
	.bot_E6END(Tile_X8Y6_E6BEG[11:0]),
	.bot_W1END(Tile_X10Y6_W1BEG[3:0]),
	.bot_W2MID(Tile_X10Y6_W2BEG[7:0]),
	.bot_W2END(Tile_X10Y6_W2BEGb[7:0]),
	.bot_WW4END(Tile_X10Y6_WW4BEG[15:0]),
	.bot_W6END(Tile_X10Y6_W6BEG[11:0]),
	.bot_E1BEG(Tile_X9Y6_E1BEG[3:0]),
	.bot_E2BEG(Tile_X9Y6_E2BEG[7:0]),
	.bot_E2BEGb(Tile_X9Y6_E2BEGb[7:0]),
	.bot_EE4BEG(Tile_X9Y6_EE4BEG[15:0]),
	.bot_E6BEG(Tile_X9Y6_E6BEG[11:0]),
	.bot_S1BEG(Tile_X9Y6_S1BEG[3:0]),
	.bot_S2BEG(Tile_X9Y6_S2BEG[7:0]),
	.bot_S2BEGb(Tile_X9Y6_S2BEGb[7:0]),
	.bot_S4BEG(Tile_X9Y6_S4BEG[15:0]),
	.bot_SS4BEG(Tile_X9Y6_SS4BEG[15:0]),
	.bot_W1BEG(Tile_X9Y6_W1BEG[3:0]),
	.bot_W2BEG(Tile_X9Y6_W2BEG[7:0]),
	.bot_W2BEGb(Tile_X9Y6_W2BEGb[7:0]),
	.bot_WW4BEG(Tile_X9Y6_WW4BEG[15:0]),
	.bot_W6BEG(Tile_X9Y6_W6BEG[11:0]),
	.UserCLK(Tile_X9Y7_UserCLKo),
	.bot_FrameData(Tile_X8Y6_FrameData_O),
	.bot_FrameData_O(Tile_X9Y6_FrameData_O),
	.FrameStrobe(Tile_X9Y7_FrameStrobe_O)
	);

	DSP Tile_X5Y7_X5Y8_DSP_tile (
	.top_E1END(Tile_X4Y7_E1BEG[3:0]),
	.top_E2MID(Tile_X4Y7_E2BEG[7:0]),
	.top_E2END(Tile_X4Y7_E2BEGb[7:0]),
	.top_EE4END(Tile_X4Y7_EE4BEG[15:0]),
	.top_E6END(Tile_X4Y7_E6BEG[11:0]),
	.top_S1END(Tile_X5Y6_S1BEG[3:0]),
	.top_S2MID(Tile_X5Y6_S2BEG[7:0]),
	.top_S2END(Tile_X5Y6_S2BEGb[7:0]),
	.top_S4END(Tile_X5Y6_S4BEG[15:0]),
	.top_SS4END(Tile_X5Y6_SS4BEG[15:0]),
	.top_W1END(Tile_X6Y7_W1BEG[3:0]),
	.top_W2MID(Tile_X6Y7_W2BEG[7:0]),
	.top_W2END(Tile_X6Y7_W2BEGb[7:0]),
	.top_WW4END(Tile_X6Y7_WW4BEG[15:0]),
	.top_W6END(Tile_X6Y7_W6BEG[11:0]),
	.top_N1BEG(Tile_X5Y7_N1BEG[3:0]),
	.top_N2BEG(Tile_X5Y7_N2BEG[7:0]),
	.top_N2BEGb(Tile_X5Y7_N2BEGb[7:0]),
	.top_N4BEG(Tile_X5Y7_N4BEG[15:0]),
	.top_NN4BEG(Tile_X5Y7_NN4BEG[15:0]),
	.top_E1BEG(Tile_X5Y7_E1BEG[3:0]),
	.top_E2BEG(Tile_X5Y7_E2BEG[7:0]),
	.top_E2BEGb(Tile_X5Y7_E2BEGb[7:0]),
	.top_EE4BEG(Tile_X5Y7_EE4BEG[15:0]),
	.top_E6BEG(Tile_X5Y7_E6BEG[11:0]),
	.top_W1BEG(Tile_X5Y7_W1BEG[3:0]),
	.top_W2BEG(Tile_X5Y7_W2BEG[7:0]),
	.top_W2BEGb(Tile_X5Y7_W2BEGb[7:0]),
	.top_WW4BEG(Tile_X5Y7_WW4BEG[15:0]),
	.top_W6BEG(Tile_X5Y7_W6BEG[11:0]),
	.top_FrameData(Tile_X4Y7_FrameData_O),
	.top_FrameData_O(Tile_X5Y7_FrameData_O),
	.FrameStrobe_O(Tile_X5Y7_FrameStrobe_O),
	.UserCLKo(Tile_X5Y7_UserCLKo),
	.bot_N1END(Tile_X5Y9_N1BEG[3:0]),
	.bot_N2MID(Tile_X5Y9_N2BEG[7:0]),
	.bot_N2END(Tile_X5Y9_N2BEGb[7:0]),
	.bot_N4END(Tile_X5Y9_N4BEG[15:0]),
	.bot_NN4END(Tile_X5Y9_NN4BEG[15:0]),
	.bot_E1END(Tile_X4Y8_E1BEG[3:0]),
	.bot_E2MID(Tile_X4Y8_E2BEG[7:0]),
	.bot_E2END(Tile_X4Y8_E2BEGb[7:0]),
	.bot_EE4END(Tile_X4Y8_EE4BEG[15:0]),
	.bot_E6END(Tile_X4Y8_E6BEG[11:0]),
	.bot_W1END(Tile_X6Y8_W1BEG[3:0]),
	.bot_W2MID(Tile_X6Y8_W2BEG[7:0]),
	.bot_W2END(Tile_X6Y8_W2BEGb[7:0]),
	.bot_WW4END(Tile_X6Y8_WW4BEG[15:0]),
	.bot_W6END(Tile_X6Y8_W6BEG[11:0]),
	.bot_E1BEG(Tile_X5Y8_E1BEG[3:0]),
	.bot_E2BEG(Tile_X5Y8_E2BEG[7:0]),
	.bot_E2BEGb(Tile_X5Y8_E2BEGb[7:0]),
	.bot_EE4BEG(Tile_X5Y8_EE4BEG[15:0]),
	.bot_E6BEG(Tile_X5Y8_E6BEG[11:0]),
	.bot_S1BEG(Tile_X5Y8_S1BEG[3:0]),
	.bot_S2BEG(Tile_X5Y8_S2BEG[7:0]),
	.bot_S2BEGb(Tile_X5Y8_S2BEGb[7:0]),
	.bot_S4BEG(Tile_X5Y8_S4BEG[15:0]),
	.bot_SS4BEG(Tile_X5Y8_SS4BEG[15:0]),
	.bot_W1BEG(Tile_X5Y8_W1BEG[3:0]),
	.bot_W2BEG(Tile_X5Y8_W2BEG[7:0]),
	.bot_W2BEGb(Tile_X5Y8_W2BEGb[7:0]),
	.bot_WW4BEG(Tile_X5Y8_WW4BEG[15:0]),
	.bot_W6BEG(Tile_X5Y8_W6BEG[11:0]),
	.UserCLK(Tile_X5Y9_UserCLKo),
	.bot_FrameData(Tile_X4Y8_FrameData_O),
	.bot_FrameData_O(Tile_X5Y8_FrameData_O),
	.FrameStrobe(Tile_X5Y9_FrameStrobe_O)
	);

	DSP Tile_X9Y7_X9Y8_DSP_tile (
	.top_E1END(Tile_X8Y7_E1BEG[3:0]),
	.top_E2MID(Tile_X8Y7_E2BEG[7:0]),
	.top_E2END(Tile_X8Y7_E2BEGb[7:0]),
	.top_EE4END(Tile_X8Y7_EE4BEG[15:0]),
	.top_E6END(Tile_X8Y7_E6BEG[11:0]),
	.top_S1END(Tile_X9Y6_S1BEG[3:0]),
	.top_S2MID(Tile_X9Y6_S2BEG[7:0]),
	.top_S2END(Tile_X9Y6_S2BEGb[7:0]),
	.top_S4END(Tile_X9Y6_S4BEG[15:0]),
	.top_SS4END(Tile_X9Y6_SS4BEG[15:0]),
	.top_W1END(Tile_X10Y7_W1BEG[3:0]),
	.top_W2MID(Tile_X10Y7_W2BEG[7:0]),
	.top_W2END(Tile_X10Y7_W2BEGb[7:0]),
	.top_WW4END(Tile_X10Y7_WW4BEG[15:0]),
	.top_W6END(Tile_X10Y7_W6BEG[11:0]),
	.top_N1BEG(Tile_X9Y7_N1BEG[3:0]),
	.top_N2BEG(Tile_X9Y7_N2BEG[7:0]),
	.top_N2BEGb(Tile_X9Y7_N2BEGb[7:0]),
	.top_N4BEG(Tile_X9Y7_N4BEG[15:0]),
	.top_NN4BEG(Tile_X9Y7_NN4BEG[15:0]),
	.top_E1BEG(Tile_X9Y7_E1BEG[3:0]),
	.top_E2BEG(Tile_X9Y7_E2BEG[7:0]),
	.top_E2BEGb(Tile_X9Y7_E2BEGb[7:0]),
	.top_EE4BEG(Tile_X9Y7_EE4BEG[15:0]),
	.top_E6BEG(Tile_X9Y7_E6BEG[11:0]),
	.top_W1BEG(Tile_X9Y7_W1BEG[3:0]),
	.top_W2BEG(Tile_X9Y7_W2BEG[7:0]),
	.top_W2BEGb(Tile_X9Y7_W2BEGb[7:0]),
	.top_WW4BEG(Tile_X9Y7_WW4BEG[15:0]),
	.top_W6BEG(Tile_X9Y7_W6BEG[11:0]),
	.top_FrameData(Tile_X8Y7_FrameData_O),
	.top_FrameData_O(Tile_X9Y7_FrameData_O),
	.FrameStrobe_O(Tile_X9Y7_FrameStrobe_O),
	.UserCLKo(Tile_X9Y7_UserCLKo),
	.bot_N1END(Tile_X9Y9_N1BEG[3:0]),
	.bot_N2MID(Tile_X9Y9_N2BEG[7:0]),
	.bot_N2END(Tile_X9Y9_N2BEGb[7:0]),
	.bot_N4END(Tile_X9Y9_N4BEG[15:0]),
	.bot_NN4END(Tile_X9Y9_NN4BEG[15:0]),
	.bot_E1END(Tile_X8Y8_E1BEG[3:0]),
	.bot_E2MID(Tile_X8Y8_E2BEG[7:0]),
	.bot_E2END(Tile_X8Y8_E2BEGb[7:0]),
	.bot_EE4END(Tile_X8Y8_EE4BEG[15:0]),
	.bot_E6END(Tile_X8Y8_E6BEG[11:0]),
	.bot_W1END(Tile_X10Y8_W1BEG[3:0]),
	.bot_W2MID(Tile_X10Y8_W2BEG[7:0]),
	.bot_W2END(Tile_X10Y8_W2BEGb[7:0]),
	.bot_WW4END(Tile_X10Y8_WW4BEG[15:0]),
	.bot_W6END(Tile_X10Y8_W6BEG[11:0]),
	.bot_E1BEG(Tile_X9Y8_E1BEG[3:0]),
	.bot_E2BEG(Tile_X9Y8_E2BEG[7:0]),
	.bot_E2BEGb(Tile_X9Y8_E2BEGb[7:0]),
	.bot_EE4BEG(Tile_X9Y8_EE4BEG[15:0]),
	.bot_E6BEG(Tile_X9Y8_E6BEG[11:0]),
	.bot_S1BEG(Tile_X9Y8_S1BEG[3:0]),
	.bot_S2BEG(Tile_X9Y8_S2BEG[7:0]),
	.bot_S2BEGb(Tile_X9Y8_S2BEGb[7:0]),
	.bot_S4BEG(Tile_X9Y8_S4BEG[15:0]),
	.bot_SS4BEG(Tile_X9Y8_SS4BEG[15:0]),
	.bot_W1BEG(Tile_X9Y8_W1BEG[3:0]),
	.bot_W2BEG(Tile_X9Y8_W2BEG[7:0]),
	.bot_W2BEGb(Tile_X9Y8_W2BEGb[7:0]),
	.bot_WW4BEG(Tile_X9Y8_WW4BEG[15:0]),
	.bot_W6BEG(Tile_X9Y8_W6BEG[11:0]),
	.UserCLK(Tile_X9Y9_UserCLKo),
	.bot_FrameData(Tile_X8Y8_FrameData_O),
	.bot_FrameData_O(Tile_X9Y8_FrameData_O),
	.FrameStrobe(Tile_X9Y9_FrameStrobe_O)
	);

	DSP Tile_X5Y9_X5Y10_DSP_tile (
	.top_E1END(Tile_X4Y9_E1BEG[3:0]),
	.top_E2MID(Tile_X4Y9_E2BEG[7:0]),
	.top_E2END(Tile_X4Y9_E2BEGb[7:0]),
	.top_EE4END(Tile_X4Y9_EE4BEG[15:0]),
	.top_E6END(Tile_X4Y9_E6BEG[11:0]),
	.top_S1END(Tile_X5Y8_S1BEG[3:0]),
	.top_S2MID(Tile_X5Y8_S2BEG[7:0]),
	.top_S2END(Tile_X5Y8_S2BEGb[7:0]),
	.top_S4END(Tile_X5Y8_S4BEG[15:0]),
	.top_SS4END(Tile_X5Y8_SS4BEG[15:0]),
	.top_W1END(Tile_X6Y9_W1BEG[3:0]),
	.top_W2MID(Tile_X6Y9_W2BEG[7:0]),
	.top_W2END(Tile_X6Y9_W2BEGb[7:0]),
	.top_WW4END(Tile_X6Y9_WW4BEG[15:0]),
	.top_W6END(Tile_X6Y9_W6BEG[11:0]),
	.top_N1BEG(Tile_X5Y9_N1BEG[3:0]),
	.top_N2BEG(Tile_X5Y9_N2BEG[7:0]),
	.top_N2BEGb(Tile_X5Y9_N2BEGb[7:0]),
	.top_N4BEG(Tile_X5Y9_N4BEG[15:0]),
	.top_NN4BEG(Tile_X5Y9_NN4BEG[15:0]),
	.top_E1BEG(Tile_X5Y9_E1BEG[3:0]),
	.top_E2BEG(Tile_X5Y9_E2BEG[7:0]),
	.top_E2BEGb(Tile_X5Y9_E2BEGb[7:0]),
	.top_EE4BEG(Tile_X5Y9_EE4BEG[15:0]),
	.top_E6BEG(Tile_X5Y9_E6BEG[11:0]),
	.top_W1BEG(Tile_X5Y9_W1BEG[3:0]),
	.top_W2BEG(Tile_X5Y9_W2BEG[7:0]),
	.top_W2BEGb(Tile_X5Y9_W2BEGb[7:0]),
	.top_WW4BEG(Tile_X5Y9_WW4BEG[15:0]),
	.top_W6BEG(Tile_X5Y9_W6BEG[11:0]),
	.top_FrameData(Tile_X4Y9_FrameData_O),
	.top_FrameData_O(Tile_X5Y9_FrameData_O),
	.FrameStrobe_O(Tile_X5Y9_FrameStrobe_O),
	.UserCLKo(Tile_X5Y9_UserCLKo),
	.bot_N1END(Tile_X5Y11_N1BEG[3:0]),
	.bot_N2MID(Tile_X5Y11_N2BEG[7:0]),
	.bot_N2END(Tile_X5Y11_N2BEGb[7:0]),
	.bot_N4END(Tile_X5Y11_N4BEG[15:0]),
	.bot_NN4END(Tile_X5Y11_NN4BEG[15:0]),
	.bot_E1END(Tile_X4Y10_E1BEG[3:0]),
	.bot_E2MID(Tile_X4Y10_E2BEG[7:0]),
	.bot_E2END(Tile_X4Y10_E2BEGb[7:0]),
	.bot_EE4END(Tile_X4Y10_EE4BEG[15:0]),
	.bot_E6END(Tile_X4Y10_E6BEG[11:0]),
	.bot_W1END(Tile_X6Y10_W1BEG[3:0]),
	.bot_W2MID(Tile_X6Y10_W2BEG[7:0]),
	.bot_W2END(Tile_X6Y10_W2BEGb[7:0]),
	.bot_WW4END(Tile_X6Y10_WW4BEG[15:0]),
	.bot_W6END(Tile_X6Y10_W6BEG[11:0]),
	.bot_E1BEG(Tile_X5Y10_E1BEG[3:0]),
	.bot_E2BEG(Tile_X5Y10_E2BEG[7:0]),
	.bot_E2BEGb(Tile_X5Y10_E2BEGb[7:0]),
	.bot_EE4BEG(Tile_X5Y10_EE4BEG[15:0]),
	.bot_E6BEG(Tile_X5Y10_E6BEG[11:0]),
	.bot_S1BEG(Tile_X5Y10_S1BEG[3:0]),
	.bot_S2BEG(Tile_X5Y10_S2BEG[7:0]),
	.bot_S2BEGb(Tile_X5Y10_S2BEGb[7:0]),
	.bot_S4BEG(Tile_X5Y10_S4BEG[15:0]),
	.bot_SS4BEG(Tile_X5Y10_SS4BEG[15:0]),
	.bot_W1BEG(Tile_X5Y10_W1BEG[3:0]),
	.bot_W2BEG(Tile_X5Y10_W2BEG[7:0]),
	.bot_W2BEGb(Tile_X5Y10_W2BEGb[7:0]),
	.bot_WW4BEG(Tile_X5Y10_WW4BEG[15:0]),
	.bot_W6BEG(Tile_X5Y10_W6BEG[11:0]),
	.UserCLK(Tile_X5Y11_UserCLKo),
	.bot_FrameData(Tile_X4Y10_FrameData_O),
	.bot_FrameData_O(Tile_X5Y10_FrameData_O),
	.FrameStrobe(Tile_X5Y11_FrameStrobe_O)
	);

	DSP Tile_X9Y9_X9Y10_DSP_tile (
	.top_E1END(Tile_X8Y9_E1BEG[3:0]),
	.top_E2MID(Tile_X8Y9_E2BEG[7:0]),
	.top_E2END(Tile_X8Y9_E2BEGb[7:0]),
	.top_EE4END(Tile_X8Y9_EE4BEG[15:0]),
	.top_E6END(Tile_X8Y9_E6BEG[11:0]),
	.top_S1END(Tile_X9Y8_S1BEG[3:0]),
	.top_S2MID(Tile_X9Y8_S2BEG[7:0]),
	.top_S2END(Tile_X9Y8_S2BEGb[7:0]),
	.top_S4END(Tile_X9Y8_S4BEG[15:0]),
	.top_SS4END(Tile_X9Y8_SS4BEG[15:0]),
	.top_W1END(Tile_X10Y9_W1BEG[3:0]),
	.top_W2MID(Tile_X10Y9_W2BEG[7:0]),
	.top_W2END(Tile_X10Y9_W2BEGb[7:0]),
	.top_WW4END(Tile_X10Y9_WW4BEG[15:0]),
	.top_W6END(Tile_X10Y9_W6BEG[11:0]),
	.top_N1BEG(Tile_X9Y9_N1BEG[3:0]),
	.top_N2BEG(Tile_X9Y9_N2BEG[7:0]),
	.top_N2BEGb(Tile_X9Y9_N2BEGb[7:0]),
	.top_N4BEG(Tile_X9Y9_N4BEG[15:0]),
	.top_NN4BEG(Tile_X9Y9_NN4BEG[15:0]),
	.top_E1BEG(Tile_X9Y9_E1BEG[3:0]),
	.top_E2BEG(Tile_X9Y9_E2BEG[7:0]),
	.top_E2BEGb(Tile_X9Y9_E2BEGb[7:0]),
	.top_EE4BEG(Tile_X9Y9_EE4BEG[15:0]),
	.top_E6BEG(Tile_X9Y9_E6BEG[11:0]),
	.top_W1BEG(Tile_X9Y9_W1BEG[3:0]),
	.top_W2BEG(Tile_X9Y9_W2BEG[7:0]),
	.top_W2BEGb(Tile_X9Y9_W2BEGb[7:0]),
	.top_WW4BEG(Tile_X9Y9_WW4BEG[15:0]),
	.top_W6BEG(Tile_X9Y9_W6BEG[11:0]),
	.top_FrameData(Tile_X8Y9_FrameData_O),
	.top_FrameData_O(Tile_X9Y9_FrameData_O),
	.FrameStrobe_O(Tile_X9Y9_FrameStrobe_O),
	.UserCLKo(Tile_X9Y9_UserCLKo),
	.bot_N1END(Tile_X9Y11_N1BEG[3:0]),
	.bot_N2MID(Tile_X9Y11_N2BEG[7:0]),
	.bot_N2END(Tile_X9Y11_N2BEGb[7:0]),
	.bot_N4END(Tile_X9Y11_N4BEG[15:0]),
	.bot_NN4END(Tile_X9Y11_NN4BEG[15:0]),
	.bot_E1END(Tile_X8Y10_E1BEG[3:0]),
	.bot_E2MID(Tile_X8Y10_E2BEG[7:0]),
	.bot_E2END(Tile_X8Y10_E2BEGb[7:0]),
	.bot_EE4END(Tile_X8Y10_EE4BEG[15:0]),
	.bot_E6END(Tile_X8Y10_E6BEG[11:0]),
	.bot_W1END(Tile_X10Y10_W1BEG[3:0]),
	.bot_W2MID(Tile_X10Y10_W2BEG[7:0]),
	.bot_W2END(Tile_X10Y10_W2BEGb[7:0]),
	.bot_WW4END(Tile_X10Y10_WW4BEG[15:0]),
	.bot_W6END(Tile_X10Y10_W6BEG[11:0]),
	.bot_E1BEG(Tile_X9Y10_E1BEG[3:0]),
	.bot_E2BEG(Tile_X9Y10_E2BEG[7:0]),
	.bot_E2BEGb(Tile_X9Y10_E2BEGb[7:0]),
	.bot_EE4BEG(Tile_X9Y10_EE4BEG[15:0]),
	.bot_E6BEG(Tile_X9Y10_E6BEG[11:0]),
	.bot_S1BEG(Tile_X9Y10_S1BEG[3:0]),
	.bot_S2BEG(Tile_X9Y10_S2BEG[7:0]),
	.bot_S2BEGb(Tile_X9Y10_S2BEGb[7:0]),
	.bot_S4BEG(Tile_X9Y10_S4BEG[15:0]),
	.bot_SS4BEG(Tile_X9Y10_SS4BEG[15:0]),
	.bot_W1BEG(Tile_X9Y10_W1BEG[3:0]),
	.bot_W2BEG(Tile_X9Y10_W2BEG[7:0]),
	.bot_W2BEGb(Tile_X9Y10_W2BEGb[7:0]),
	.bot_WW4BEG(Tile_X9Y10_WW4BEG[15:0]),
	.bot_W6BEG(Tile_X9Y10_W6BEG[11:0]),
	.UserCLK(Tile_X9Y11_UserCLKo),
	.bot_FrameData(Tile_X8Y10_FrameData_O),
	.bot_FrameData_O(Tile_X9Y10_FrameData_O),
	.FrameStrobe(Tile_X9Y11_FrameStrobe_O)
	);

	DSP Tile_X5Y11_X5Y12_DSP_tile (
	.top_E1END(Tile_X4Y11_E1BEG[3:0]),
	.top_E2MID(Tile_X4Y11_E2BEG[7:0]),
	.top_E2END(Tile_X4Y11_E2BEGb[7:0]),
	.top_EE4END(Tile_X4Y11_EE4BEG[15:0]),
	.top_E6END(Tile_X4Y11_E6BEG[11:0]),
	.top_S1END(Tile_X5Y10_S1BEG[3:0]),
	.top_S2MID(Tile_X5Y10_S2BEG[7:0]),
	.top_S2END(Tile_X5Y10_S2BEGb[7:0]),
	.top_S4END(Tile_X5Y10_S4BEG[15:0]),
	.top_SS4END(Tile_X5Y10_SS4BEG[15:0]),
	.top_W1END(Tile_X6Y11_W1BEG[3:0]),
	.top_W2MID(Tile_X6Y11_W2BEG[7:0]),
	.top_W2END(Tile_X6Y11_W2BEGb[7:0]),
	.top_WW4END(Tile_X6Y11_WW4BEG[15:0]),
	.top_W6END(Tile_X6Y11_W6BEG[11:0]),
	.top_N1BEG(Tile_X5Y11_N1BEG[3:0]),
	.top_N2BEG(Tile_X5Y11_N2BEG[7:0]),
	.top_N2BEGb(Tile_X5Y11_N2BEGb[7:0]),
	.top_N4BEG(Tile_X5Y11_N4BEG[15:0]),
	.top_NN4BEG(Tile_X5Y11_NN4BEG[15:0]),
	.top_E1BEG(Tile_X5Y11_E1BEG[3:0]),
	.top_E2BEG(Tile_X5Y11_E2BEG[7:0]),
	.top_E2BEGb(Tile_X5Y11_E2BEGb[7:0]),
	.top_EE4BEG(Tile_X5Y11_EE4BEG[15:0]),
	.top_E6BEG(Tile_X5Y11_E6BEG[11:0]),
	.top_W1BEG(Tile_X5Y11_W1BEG[3:0]),
	.top_W2BEG(Tile_X5Y11_W2BEG[7:0]),
	.top_W2BEGb(Tile_X5Y11_W2BEGb[7:0]),
	.top_WW4BEG(Tile_X5Y11_WW4BEG[15:0]),
	.top_W6BEG(Tile_X5Y11_W6BEG[11:0]),
	.top_FrameData(Tile_X4Y11_FrameData_O),
	.top_FrameData_O(Tile_X5Y11_FrameData_O),
	.FrameStrobe_O(Tile_X5Y11_FrameStrobe_O),
	.UserCLKo(Tile_X5Y11_UserCLKo),
	.bot_N1END(Tile_X5Y13_N1BEG[3:0]),
	.bot_N2MID(Tile_X5Y13_N2BEG[7:0]),
	.bot_N2END(Tile_X5Y13_N2BEGb[7:0]),
	.bot_N4END(Tile_X5Y13_N4BEG[15:0]),
	.bot_NN4END(Tile_X5Y13_NN4BEG[15:0]),
	.bot_E1END(Tile_X4Y12_E1BEG[3:0]),
	.bot_E2MID(Tile_X4Y12_E2BEG[7:0]),
	.bot_E2END(Tile_X4Y12_E2BEGb[7:0]),
	.bot_EE4END(Tile_X4Y12_EE4BEG[15:0]),
	.bot_E6END(Tile_X4Y12_E6BEG[11:0]),
	.bot_W1END(Tile_X6Y12_W1BEG[3:0]),
	.bot_W2MID(Tile_X6Y12_W2BEG[7:0]),
	.bot_W2END(Tile_X6Y12_W2BEGb[7:0]),
	.bot_WW4END(Tile_X6Y12_WW4BEG[15:0]),
	.bot_W6END(Tile_X6Y12_W6BEG[11:0]),
	.bot_E1BEG(Tile_X5Y12_E1BEG[3:0]),
	.bot_E2BEG(Tile_X5Y12_E2BEG[7:0]),
	.bot_E2BEGb(Tile_X5Y12_E2BEGb[7:0]),
	.bot_EE4BEG(Tile_X5Y12_EE4BEG[15:0]),
	.bot_E6BEG(Tile_X5Y12_E6BEG[11:0]),
	.bot_S1BEG(Tile_X5Y12_S1BEG[3:0]),
	.bot_S2BEG(Tile_X5Y12_S2BEG[7:0]),
	.bot_S2BEGb(Tile_X5Y12_S2BEGb[7:0]),
	.bot_S4BEG(Tile_X5Y12_S4BEG[15:0]),
	.bot_SS4BEG(Tile_X5Y12_SS4BEG[15:0]),
	.bot_W1BEG(Tile_X5Y12_W1BEG[3:0]),
	.bot_W2BEG(Tile_X5Y12_W2BEG[7:0]),
	.bot_W2BEGb(Tile_X5Y12_W2BEGb[7:0]),
	.bot_WW4BEG(Tile_X5Y12_WW4BEG[15:0]),
	.bot_W6BEG(Tile_X5Y12_W6BEG[11:0]),
	.UserCLK(Tile_X5Y13_UserCLKo),
	.bot_FrameData(Tile_X4Y12_FrameData_O),
	.bot_FrameData_O(Tile_X5Y12_FrameData_O),
	.FrameStrobe(Tile_X5Y13_FrameStrobe_O)
	);

	DSP Tile_X9Y11_X9Y12_DSP_tile (
	.top_E1END(Tile_X8Y11_E1BEG[3:0]),
	.top_E2MID(Tile_X8Y11_E2BEG[7:0]),
	.top_E2END(Tile_X8Y11_E2BEGb[7:0]),
	.top_EE4END(Tile_X8Y11_EE4BEG[15:0]),
	.top_E6END(Tile_X8Y11_E6BEG[11:0]),
	.top_S1END(Tile_X9Y10_S1BEG[3:0]),
	.top_S2MID(Tile_X9Y10_S2BEG[7:0]),
	.top_S2END(Tile_X9Y10_S2BEGb[7:0]),
	.top_S4END(Tile_X9Y10_S4BEG[15:0]),
	.top_SS4END(Tile_X9Y10_SS4BEG[15:0]),
	.top_W1END(Tile_X10Y11_W1BEG[3:0]),
	.top_W2MID(Tile_X10Y11_W2BEG[7:0]),
	.top_W2END(Tile_X10Y11_W2BEGb[7:0]),
	.top_WW4END(Tile_X10Y11_WW4BEG[15:0]),
	.top_W6END(Tile_X10Y11_W6BEG[11:0]),
	.top_N1BEG(Tile_X9Y11_N1BEG[3:0]),
	.top_N2BEG(Tile_X9Y11_N2BEG[7:0]),
	.top_N2BEGb(Tile_X9Y11_N2BEGb[7:0]),
	.top_N4BEG(Tile_X9Y11_N4BEG[15:0]),
	.top_NN4BEG(Tile_X9Y11_NN4BEG[15:0]),
	.top_E1BEG(Tile_X9Y11_E1BEG[3:0]),
	.top_E2BEG(Tile_X9Y11_E2BEG[7:0]),
	.top_E2BEGb(Tile_X9Y11_E2BEGb[7:0]),
	.top_EE4BEG(Tile_X9Y11_EE4BEG[15:0]),
	.top_E6BEG(Tile_X9Y11_E6BEG[11:0]),
	.top_W1BEG(Tile_X9Y11_W1BEG[3:0]),
	.top_W2BEG(Tile_X9Y11_W2BEG[7:0]),
	.top_W2BEGb(Tile_X9Y11_W2BEGb[7:0]),
	.top_WW4BEG(Tile_X9Y11_WW4BEG[15:0]),
	.top_W6BEG(Tile_X9Y11_W6BEG[11:0]),
	.top_FrameData(Tile_X8Y11_FrameData_O),
	.top_FrameData_O(Tile_X9Y11_FrameData_O),
	.FrameStrobe_O(Tile_X9Y11_FrameStrobe_O),
	.UserCLKo(Tile_X9Y11_UserCLKo),
	.bot_N1END(Tile_X9Y13_N1BEG[3:0]),
	.bot_N2MID(Tile_X9Y13_N2BEG[7:0]),
	.bot_N2END(Tile_X9Y13_N2BEGb[7:0]),
	.bot_N4END(Tile_X9Y13_N4BEG[15:0]),
	.bot_NN4END(Tile_X9Y13_NN4BEG[15:0]),
	.bot_E1END(Tile_X8Y12_E1BEG[3:0]),
	.bot_E2MID(Tile_X8Y12_E2BEG[7:0]),
	.bot_E2END(Tile_X8Y12_E2BEGb[7:0]),
	.bot_EE4END(Tile_X8Y12_EE4BEG[15:0]),
	.bot_E6END(Tile_X8Y12_E6BEG[11:0]),
	.bot_W1END(Tile_X10Y12_W1BEG[3:0]),
	.bot_W2MID(Tile_X10Y12_W2BEG[7:0]),
	.bot_W2END(Tile_X10Y12_W2BEGb[7:0]),
	.bot_WW4END(Tile_X10Y12_WW4BEG[15:0]),
	.bot_W6END(Tile_X10Y12_W6BEG[11:0]),
	.bot_E1BEG(Tile_X9Y12_E1BEG[3:0]),
	.bot_E2BEG(Tile_X9Y12_E2BEG[7:0]),
	.bot_E2BEGb(Tile_X9Y12_E2BEGb[7:0]),
	.bot_EE4BEG(Tile_X9Y12_EE4BEG[15:0]),
	.bot_E6BEG(Tile_X9Y12_E6BEG[11:0]),
	.bot_S1BEG(Tile_X9Y12_S1BEG[3:0]),
	.bot_S2BEG(Tile_X9Y12_S2BEG[7:0]),
	.bot_S2BEGb(Tile_X9Y12_S2BEGb[7:0]),
	.bot_S4BEG(Tile_X9Y12_S4BEG[15:0]),
	.bot_SS4BEG(Tile_X9Y12_SS4BEG[15:0]),
	.bot_W1BEG(Tile_X9Y12_W1BEG[3:0]),
	.bot_W2BEG(Tile_X9Y12_W2BEG[7:0]),
	.bot_W2BEGb(Tile_X9Y12_W2BEGb[7:0]),
	.bot_WW4BEG(Tile_X9Y12_WW4BEG[15:0]),
	.bot_W6BEG(Tile_X9Y12_W6BEG[11:0]),
	.UserCLK(Tile_X9Y13_UserCLKo),
	.bot_FrameData(Tile_X8Y12_FrameData_O),
	.bot_FrameData_O(Tile_X9Y12_FrameData_O),
	.FrameStrobe(Tile_X9Y13_FrameStrobe_O)
	);

endmodule
