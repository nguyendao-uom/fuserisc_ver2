magic
tech sky130A
magscale 1 2
timestamp 1637968891
<< locali >>
rect 582389 677535 582423 697153
rect 582389 648567 582423 670701
rect 582481 662371 582515 683825
rect 582389 633403 582423 643977
rect 582389 618239 582423 630785
rect 582389 604435 582423 617457
rect 582389 575467 582423 577609
rect 582389 560235 582423 564281
rect 582389 537863 582423 543745
rect 582389 524535 582423 529941
rect 582389 511343 582423 514913
rect 582389 484687 582423 500973
rect 582481 471495 582515 485809
rect 582573 458167 582607 470781
rect 582389 431647 582423 456773
rect 582481 418319 582515 442017
rect 582389 378471 582423 412777
rect 582573 404991 582607 426445
rect 582389 325295 582423 368509
rect 582481 365143 582515 397477
rect 582573 351951 582607 383673
rect 582389 258927 582423 310505
rect 582481 272255 582515 324309
rect 582573 298775 582607 339473
rect 582665 312103 582699 353277
rect 582389 205751 582423 251209
rect 582481 219079 582515 266373
rect 582573 245599 582607 295341
rect 582665 232407 582699 280177
rect 582389 126055 582423 162877
rect 582481 139383 582515 178041
rect 582573 152711 582607 193205
rect 582665 179231 582699 222173
rect 582757 192559 582791 235977
rect 582849 165903 582883 207009
rect 582389 86207 582423 118677
rect 582481 99535 582515 133909
rect 582573 112863 582607 149073
rect 582389 46359 582423 75905
rect 582481 59687 582515 89709
rect 582573 73015 582607 104873
rect 582573 33099 582607 60741
rect 83565 27251 83599 27421
rect 582481 6647 582515 31773
rect 582665 19839 582699 46121
<< viali >>
rect 582389 697153 582423 697187
rect 582389 677501 582423 677535
rect 582481 683825 582515 683859
rect 582389 670701 582423 670735
rect 582481 662337 582515 662371
rect 582389 648533 582423 648567
rect 582389 643977 582423 644011
rect 582389 633369 582423 633403
rect 582389 630785 582423 630819
rect 582389 618205 582423 618239
rect 582389 617457 582423 617491
rect 582389 604401 582423 604435
rect 582389 577609 582423 577643
rect 582389 575433 582423 575467
rect 582389 564281 582423 564315
rect 582389 560201 582423 560235
rect 582389 543745 582423 543779
rect 582389 537829 582423 537863
rect 582389 529941 582423 529975
rect 582389 524501 582423 524535
rect 582389 514913 582423 514947
rect 582389 511309 582423 511343
rect 582389 500973 582423 501007
rect 582389 484653 582423 484687
rect 582481 485809 582515 485843
rect 582481 471461 582515 471495
rect 582573 470781 582607 470815
rect 582573 458133 582607 458167
rect 582389 456773 582423 456807
rect 582389 431613 582423 431647
rect 582481 442017 582515 442051
rect 582481 418285 582515 418319
rect 582573 426445 582607 426479
rect 582389 412777 582423 412811
rect 582573 404957 582607 404991
rect 582389 378437 582423 378471
rect 582481 397477 582515 397511
rect 582389 368509 582423 368543
rect 582481 365109 582515 365143
rect 582573 383673 582607 383707
rect 582573 351917 582607 351951
rect 582665 353277 582699 353311
rect 582389 325261 582423 325295
rect 582573 339473 582607 339507
rect 582481 324309 582515 324343
rect 582389 310505 582423 310539
rect 582665 312069 582699 312103
rect 582573 298741 582607 298775
rect 582481 272221 582515 272255
rect 582573 295341 582607 295375
rect 582389 258893 582423 258927
rect 582481 266373 582515 266407
rect 582389 251209 582423 251243
rect 582573 245565 582607 245599
rect 582665 280177 582699 280211
rect 582665 232373 582699 232407
rect 582757 235977 582791 236011
rect 582481 219045 582515 219079
rect 582665 222173 582699 222207
rect 582389 205717 582423 205751
rect 582573 193205 582607 193239
rect 582481 178041 582515 178075
rect 582389 162877 582423 162911
rect 582757 192525 582791 192559
rect 582849 207009 582883 207043
rect 582665 179197 582699 179231
rect 582849 165869 582883 165903
rect 582573 152677 582607 152711
rect 582481 139349 582515 139383
rect 582573 149073 582607 149107
rect 582389 126021 582423 126055
rect 582481 133909 582515 133943
rect 582389 118677 582423 118711
rect 582573 112829 582607 112863
rect 582481 99501 582515 99535
rect 582573 104873 582607 104907
rect 582389 86173 582423 86207
rect 582481 89709 582515 89743
rect 582389 75905 582423 75939
rect 582573 72981 582607 73015
rect 582481 59653 582515 59687
rect 582573 60741 582607 60775
rect 582389 46325 582423 46359
rect 582573 33065 582607 33099
rect 582665 46121 582699 46155
rect 582481 31773 582515 31807
rect 83565 27421 83599 27455
rect 83565 27217 83599 27251
rect 582665 19805 582699 19839
rect 582481 6613 582515 6647
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 364978 700476 364984 700528
rect 365036 700516 365042 700528
rect 365622 700516 365628 700528
rect 365036 700488 365628 700516
rect 365036 700476 365042 700488
rect 365622 700476 365628 700488
rect 365680 700476 365686 700528
rect 527174 700476 527180 700528
rect 527232 700516 527238 700528
rect 528462 700516 528468 700528
rect 527232 700488 528468 700516
rect 527232 700476 527238 700488
rect 528462 700476 528468 700488
rect 528520 700476 528526 700528
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 105446 700340 105452 700392
rect 105504 700380 105510 700392
rect 106182 700380 106188 700392
rect 105504 700352 106188 700380
rect 105504 700340 105510 700352
rect 106182 700340 106188 700352
rect 106240 700340 106246 700392
rect 235166 700340 235172 700392
rect 235224 700380 235230 700392
rect 235902 700380 235908 700392
rect 235224 700352 235908 700380
rect 235224 700340 235230 700352
rect 235902 700340 235908 700352
rect 235960 700340 235966 700392
rect 170306 700204 170312 700256
rect 170364 700244 170370 700256
rect 171042 700244 171048 700256
rect 170364 700216 171048 700244
rect 170364 700204 170370 700216
rect 171042 700204 171048 700216
rect 171100 700204 171106 700256
rect 397454 699932 397460 699984
rect 397512 699972 397518 699984
rect 398742 699972 398748 699984
rect 397512 699944 398748 699972
rect 397512 699932 397518 699944
rect 398742 699932 398748 699944
rect 398800 699932 398806 699984
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 300762 699700 300768 699712
rect 300176 699672 300768 699700
rect 300176 699660 300182 699672
rect 300762 699660 300768 699672
rect 300820 699660 300826 699712
rect 429838 699660 429844 699712
rect 429896 699700 429902 699712
rect 430482 699700 430488 699712
rect 429896 699672 430488 699700
rect 429896 699660 429902 699672
rect 430482 699660 430488 699672
rect 430540 699660 430546 699712
rect 462314 699660 462320 699712
rect 462372 699700 462378 699712
rect 463602 699700 463608 699712
rect 462372 699672 463608 699700
rect 462372 699660 462378 699672
rect 463602 699660 463608 699672
rect 463660 699660 463666 699712
rect 494790 699660 494796 699712
rect 494848 699700 494854 699712
rect 495342 699700 495348 699712
rect 494848 699672 495348 699700
rect 494848 699660 494854 699672
rect 495342 699660 495348 699672
rect 495400 699660 495406 699712
rect 559650 699660 559656 699712
rect 559708 699700 559714 699712
rect 560202 699700 560208 699712
rect 559708 699672 560208 699700
rect 559708 699660 559714 699672
rect 560202 699660 560208 699672
rect 560260 699660 560266 699712
rect 582374 697184 582380 697196
rect 582335 697156 582380 697184
rect 582374 697144 582380 697156
rect 582432 697144 582438 697196
rect 582466 683856 582472 683868
rect 582427 683828 582472 683856
rect 582466 683816 582472 683828
rect 582524 683816 582530 683868
rect 6086 681640 6092 681692
rect 6144 681680 6150 681692
rect 6914 681680 6920 681692
rect 6144 681652 6920 681680
rect 6144 681640 6150 681652
rect 6914 681640 6920 681652
rect 6972 681640 6978 681692
rect 24762 681640 24768 681692
rect 24820 681680 24826 681692
rect 27982 681680 27988 681692
rect 24820 681652 27988 681680
rect 24820 681640 24826 681652
rect 27982 681640 27988 681652
rect 28040 681640 28046 681692
rect 89622 681640 89628 681692
rect 89680 681680 89686 681692
rect 93946 681680 93952 681692
rect 89680 681652 93952 681680
rect 89680 681640 89686 681652
rect 93946 681640 93952 681652
rect 94004 681640 94010 681692
rect 267642 681232 267648 681284
rect 267700 681272 267706 681284
rect 270034 681272 270040 681284
rect 267700 681244 270040 681272
rect 267700 681232 267706 681244
rect 270034 681232 270040 681244
rect 270092 681232 270098 681284
rect 332502 681096 332508 681148
rect 332560 681136 332566 681148
rect 335998 681136 336004 681148
rect 332560 681108 336004 681136
rect 332560 681096 332566 681108
rect 335998 681096 336004 681108
rect 336056 681096 336062 681148
rect 41322 680960 41328 681012
rect 41380 681000 41386 681012
rect 49970 681000 49976 681012
rect 41380 680972 49976 681000
rect 41380 680960 41386 680972
rect 49970 680960 49976 680972
rect 50028 680960 50034 681012
rect 106182 680960 106188 681012
rect 106240 681000 106246 681012
rect 115934 681000 115940 681012
rect 106240 680972 115940 681000
rect 106240 680960 106246 680972
rect 115934 680960 115940 680972
rect 115992 680960 115998 681012
rect 171042 680960 171048 681012
rect 171100 681000 171106 681012
rect 181990 681000 181996 681012
rect 171100 680972 181996 681000
rect 171100 680960 171106 680972
rect 181990 680960 181996 680972
rect 182048 680960 182054 681012
rect 219342 680960 219348 681012
rect 219400 681000 219406 681012
rect 225966 681000 225972 681012
rect 219400 680972 225972 681000
rect 219400 680960 219406 680972
rect 225966 680960 225972 680972
rect 226024 680960 226030 681012
rect 235902 680960 235908 681012
rect 235960 681000 235966 681012
rect 248046 681000 248052 681012
rect 235960 680972 248052 681000
rect 235960 680960 235966 680972
rect 248046 680960 248052 680972
rect 248104 680960 248110 681012
rect 284202 680960 284208 681012
rect 284260 681000 284266 681012
rect 292022 681000 292028 681012
rect 284260 680972 292028 681000
rect 284260 680960 284266 680972
rect 292022 680960 292028 680972
rect 292080 680960 292086 681012
rect 300762 680960 300768 681012
rect 300820 681000 300826 681012
rect 314010 681000 314016 681012
rect 300820 680972 314016 681000
rect 300820 680960 300826 680972
rect 314010 680960 314016 680972
rect 314068 680960 314074 681012
rect 349062 680960 349068 681012
rect 349120 681000 349126 681012
rect 358078 681000 358084 681012
rect 349120 680972 358084 681000
rect 349120 680960 349126 680972
rect 358078 680960 358084 680972
rect 358136 680960 358142 681012
rect 365622 680960 365628 681012
rect 365680 681000 365686 681012
rect 380066 681000 380072 681012
rect 365680 680972 380072 681000
rect 365680 680960 365686 680972
rect 380066 680960 380072 680972
rect 380124 680960 380130 681012
rect 413922 680960 413928 681012
rect 413980 681000 413986 681012
rect 424042 681000 424048 681012
rect 413980 680972 424048 681000
rect 413980 680960 413986 680972
rect 424042 680960 424048 680972
rect 424100 680960 424106 681012
rect 430482 680960 430488 681012
rect 430540 681000 430546 681012
rect 446030 681000 446036 681012
rect 430540 680972 446036 681000
rect 430540 680960 430546 680972
rect 446030 680960 446036 680972
rect 446088 680960 446094 681012
rect 478782 680960 478788 681012
rect 478840 681000 478846 681012
rect 490098 681000 490104 681012
rect 478840 680972 490104 681000
rect 478840 680960 478846 680972
rect 490098 680960 490104 680972
rect 490156 680960 490162 681012
rect 495342 680960 495348 681012
rect 495400 681000 495406 681012
rect 512086 681000 512092 681012
rect 495400 680972 512092 681000
rect 495400 680960 495406 680972
rect 512086 680960 512092 680972
rect 512144 680960 512150 681012
rect 528462 680960 528468 681012
rect 528520 681000 528526 681012
rect 534074 681000 534080 681012
rect 528520 680972 534080 681000
rect 528520 680960 528526 680972
rect 534074 680960 534080 680972
rect 534132 680960 534138 681012
rect 543642 680960 543648 681012
rect 543700 681000 543706 681012
rect 556062 681000 556068 681012
rect 543700 680972 556068 681000
rect 543700 680960 543706 680972
rect 556062 680960 556068 680972
rect 556120 680960 556126 681012
rect 560202 680960 560208 681012
rect 560260 681000 560266 681012
rect 578050 681000 578056 681012
rect 560260 680972 578056 681000
rect 560260 680960 560266 680972
rect 578050 680960 578056 680972
rect 578108 680960 578114 681012
rect 202782 680892 202788 680944
rect 202840 680932 202846 680944
rect 203978 680932 203984 680944
rect 202840 680904 203984 680932
rect 202840 680892 202846 680904
rect 203978 680892 203984 680904
rect 204036 680892 204042 680944
rect 463602 680892 463608 680944
rect 463660 680932 463666 680944
rect 468110 680932 468116 680944
rect 463660 680904 468116 680932
rect 463660 680892 463666 680904
rect 468110 680892 468116 680904
rect 468168 680892 468174 680944
rect 398742 680688 398748 680740
rect 398800 680728 398806 680740
rect 402054 680728 402060 680740
rect 398800 680700 402060 680728
rect 398800 680688 398806 680700
rect 402054 680688 402060 680700
rect 402112 680688 402118 680740
rect 154482 680620 154488 680672
rect 154540 680660 154546 680672
rect 160002 680660 160008 680672
rect 154540 680632 160008 680660
rect 154540 680620 154546 680632
rect 160002 680620 160008 680632
rect 160060 680620 160066 680672
rect 582374 677532 582380 677544
rect 582335 677504 582380 677532
rect 582374 677492 582380 677504
rect 582432 677492 582438 677544
rect 582374 670732 582380 670744
rect 582335 670704 582380 670732
rect 582374 670692 582380 670704
rect 582432 670692 582438 670744
rect 582466 662368 582472 662380
rect 582427 662340 582472 662368
rect 582466 662328 582472 662340
rect 582524 662328 582530 662380
rect 106 658180 112 658232
rect 164 658220 170 658232
rect 566 658220 572 658232
rect 164 658192 572 658220
rect 164 658180 170 658192
rect 566 658180 572 658192
rect 624 658180 630 658232
rect 582374 648564 582380 648576
rect 582335 648536 582380 648564
rect 582374 648524 582380 648536
rect 582432 648524 582438 648576
rect 582374 644008 582380 644020
rect 582335 643980 582380 644008
rect 582374 643968 582380 643980
rect 582432 643968 582438 644020
rect 582374 633400 582380 633412
rect 582335 633372 582380 633400
rect 582374 633360 582380 633372
rect 582432 633360 582438 633412
rect 14 632068 20 632120
rect 72 632108 78 632120
rect 566 632108 572 632120
rect 72 632080 572 632108
rect 72 632068 78 632080
rect 566 632068 572 632080
rect 624 632068 630 632120
rect 582374 630816 582380 630828
rect 582335 630788 582380 630816
rect 582374 630776 582380 630788
rect 582432 630776 582438 630828
rect 582374 618236 582380 618248
rect 582335 618208 582380 618236
rect 582374 618196 582380 618208
rect 582432 618196 582438 618248
rect 582374 617488 582380 617500
rect 582335 617460 582380 617488
rect 582374 617448 582380 617460
rect 582432 617448 582438 617500
rect 582374 604432 582380 604444
rect 582335 604404 582380 604432
rect 582374 604392 582380 604404
rect 582432 604392 582438 604444
rect 582374 577640 582380 577652
rect 582335 577612 582380 577640
rect 582374 577600 582380 577612
rect 582432 577600 582438 577652
rect 582374 575464 582380 575476
rect 582335 575436 582380 575464
rect 582374 575424 582380 575436
rect 582432 575424 582438 575476
rect 582374 564312 582380 564324
rect 582335 564284 582380 564312
rect 582374 564272 582380 564284
rect 582432 564272 582438 564324
rect 582374 560232 582380 560244
rect 582335 560204 582380 560232
rect 582374 560192 582380 560204
rect 582432 560192 582438 560244
rect 582374 543776 582380 543788
rect 582335 543748 582380 543776
rect 582374 543736 582380 543748
rect 582432 543736 582438 543788
rect 582374 537860 582380 537872
rect 582335 537832 582380 537860
rect 582374 537820 582380 537832
rect 582432 537820 582438 537872
rect 582374 529972 582380 529984
rect 582335 529944 582380 529972
rect 582374 529932 582380 529944
rect 582432 529932 582438 529984
rect 582374 524532 582380 524544
rect 582335 524504 582380 524532
rect 582374 524492 582380 524504
rect 582432 524492 582438 524544
rect 582374 514944 582380 514956
rect 582335 514916 582380 514944
rect 582374 514904 582380 514916
rect 582432 514904 582438 514956
rect 582374 511340 582380 511352
rect 582335 511312 582380 511340
rect 582374 511300 582380 511312
rect 582432 511300 582438 511352
rect 582374 501004 582380 501016
rect 582335 500976 582380 501004
rect 582374 500964 582380 500976
rect 582432 500964 582438 501016
rect 582466 485840 582472 485852
rect 582427 485812 582472 485840
rect 582466 485800 582472 485812
rect 582524 485800 582530 485852
rect 582374 484684 582380 484696
rect 582335 484656 582380 484684
rect 582374 484644 582380 484656
rect 582432 484644 582438 484696
rect 582466 471492 582472 471504
rect 582427 471464 582472 471492
rect 582466 471452 582472 471464
rect 582524 471452 582530 471504
rect 582558 470812 582564 470824
rect 582519 470784 582564 470812
rect 582558 470772 582564 470784
rect 582616 470772 582622 470824
rect 582558 458164 582564 458176
rect 582519 458136 582564 458164
rect 582558 458124 582564 458136
rect 582616 458124 582622 458176
rect 582374 456804 582380 456816
rect 582335 456776 582380 456804
rect 582374 456764 582380 456776
rect 582432 456764 582438 456816
rect 582466 442048 582472 442060
rect 582427 442020 582472 442048
rect 582466 442008 582472 442020
rect 582524 442008 582530 442060
rect 582374 431644 582380 431656
rect 582335 431616 582380 431644
rect 582374 431604 582380 431616
rect 582432 431604 582438 431656
rect 582558 426476 582564 426488
rect 582519 426448 582564 426476
rect 582558 426436 582564 426448
rect 582616 426436 582622 426488
rect 582466 418316 582472 418328
rect 582427 418288 582472 418316
rect 582466 418276 582472 418288
rect 582524 418276 582530 418328
rect 582374 412808 582380 412820
rect 582335 412780 582380 412808
rect 582374 412768 582380 412780
rect 582432 412768 582438 412820
rect 582558 404988 582564 405000
rect 582519 404960 582564 404988
rect 582558 404948 582564 404960
rect 582616 404948 582622 405000
rect 582466 397508 582472 397520
rect 582427 397480 582472 397508
rect 582466 397468 582472 397480
rect 582524 397468 582530 397520
rect 582558 383704 582564 383716
rect 582519 383676 582564 383704
rect 582558 383664 582564 383676
rect 582616 383664 582622 383716
rect 582374 378468 582380 378480
rect 582335 378440 582380 378468
rect 582374 378428 582380 378440
rect 582432 378428 582438 378480
rect 582374 368540 582380 368552
rect 582335 368512 582380 368540
rect 582374 368500 582380 368512
rect 582432 368500 582438 368552
rect 582466 365140 582472 365152
rect 582427 365112 582472 365140
rect 582466 365100 582472 365112
rect 582524 365100 582530 365152
rect 582650 353308 582656 353320
rect 582611 353280 582656 353308
rect 582650 353268 582656 353280
rect 582708 353268 582714 353320
rect 582558 351948 582564 351960
rect 582519 351920 582564 351948
rect 582558 351908 582564 351920
rect 582616 351908 582622 351960
rect 582558 339504 582564 339516
rect 582519 339476 582564 339504
rect 582558 339464 582564 339476
rect 582616 339464 582622 339516
rect 582374 325292 582380 325304
rect 582335 325264 582380 325292
rect 582374 325252 582380 325264
rect 582432 325252 582438 325304
rect 582466 324340 582472 324352
rect 582427 324312 582472 324340
rect 582466 324300 582472 324312
rect 582524 324300 582530 324352
rect 582650 312100 582656 312112
rect 582611 312072 582656 312100
rect 582650 312060 582656 312072
rect 582708 312060 582714 312112
rect 582374 310536 582380 310548
rect 582335 310508 582380 310536
rect 582374 310496 582380 310508
rect 582432 310496 582438 310548
rect 582558 298772 582564 298784
rect 582519 298744 582564 298772
rect 582558 298732 582564 298744
rect 582616 298732 582622 298784
rect 582558 295372 582564 295384
rect 582519 295344 582564 295372
rect 582558 295332 582564 295344
rect 582616 295332 582622 295384
rect 582650 280208 582656 280220
rect 582611 280180 582656 280208
rect 582650 280168 582656 280180
rect 582708 280168 582714 280220
rect 582466 272252 582472 272264
rect 582427 272224 582472 272252
rect 582466 272212 582472 272224
rect 582524 272212 582530 272264
rect 582466 266404 582472 266416
rect 582427 266376 582472 266404
rect 582466 266364 582472 266376
rect 582524 266364 582530 266416
rect 582374 258924 582380 258936
rect 582335 258896 582380 258924
rect 582374 258884 582380 258896
rect 582432 258884 582438 258936
rect 582374 251240 582380 251252
rect 582335 251212 582380 251240
rect 582374 251200 582380 251212
rect 582432 251200 582438 251252
rect 582558 245596 582564 245608
rect 582519 245568 582564 245596
rect 582558 245556 582564 245568
rect 582616 245556 582622 245608
rect 582742 236008 582748 236020
rect 582703 235980 582748 236008
rect 582742 235968 582748 235980
rect 582800 235968 582806 236020
rect 582650 232404 582656 232416
rect 582611 232376 582656 232404
rect 582650 232364 582656 232376
rect 582708 232364 582714 232416
rect 582650 222204 582656 222216
rect 582611 222176 582656 222204
rect 582650 222164 582656 222176
rect 582708 222164 582714 222216
rect 582466 219076 582472 219088
rect 582427 219048 582472 219076
rect 582466 219036 582472 219048
rect 582524 219036 582530 219088
rect 582834 207040 582840 207052
rect 582795 207012 582840 207040
rect 582834 207000 582840 207012
rect 582892 207000 582898 207052
rect 582374 205748 582380 205760
rect 582335 205720 582380 205748
rect 582374 205708 582380 205720
rect 582432 205708 582438 205760
rect 582558 193236 582564 193248
rect 582519 193208 582564 193236
rect 582558 193196 582564 193208
rect 582616 193196 582622 193248
rect 582742 192556 582748 192568
rect 582703 192528 582748 192556
rect 582742 192516 582748 192528
rect 582800 192516 582806 192568
rect 582650 179228 582656 179240
rect 582611 179200 582656 179228
rect 582650 179188 582656 179200
rect 582708 179188 582714 179240
rect 582466 178072 582472 178084
rect 582427 178044 582472 178072
rect 582466 178032 582472 178044
rect 582524 178032 582530 178084
rect 582834 165900 582840 165912
rect 582795 165872 582840 165900
rect 582834 165860 582840 165872
rect 582892 165860 582898 165912
rect 582374 162908 582380 162920
rect 582335 162880 582380 162908
rect 582374 162868 582380 162880
rect 582432 162868 582438 162920
rect 582558 152708 582564 152720
rect 582519 152680 582564 152708
rect 582558 152668 582564 152680
rect 582616 152668 582622 152720
rect 582558 149104 582564 149116
rect 582519 149076 582564 149104
rect 582558 149064 582564 149076
rect 582616 149064 582622 149116
rect 582466 139380 582472 139392
rect 582427 139352 582472 139380
rect 582466 139340 582472 139352
rect 582524 139340 582530 139392
rect 582466 133940 582472 133952
rect 582427 133912 582472 133940
rect 582466 133900 582472 133912
rect 582524 133900 582530 133952
rect 582374 126052 582380 126064
rect 582335 126024 582380 126052
rect 582374 126012 582380 126024
rect 582432 126012 582438 126064
rect 582374 118708 582380 118720
rect 582335 118680 582380 118708
rect 582374 118668 582380 118680
rect 582432 118668 582438 118720
rect 582558 112860 582564 112872
rect 582519 112832 582564 112860
rect 582558 112820 582564 112832
rect 582616 112820 582622 112872
rect 582558 104904 582564 104916
rect 582519 104876 582564 104904
rect 582558 104864 582564 104876
rect 582616 104864 582622 104916
rect 582466 99532 582472 99544
rect 582427 99504 582472 99532
rect 582466 99492 582472 99504
rect 582524 99492 582530 99544
rect 582466 89740 582472 89752
rect 582427 89712 582472 89740
rect 582466 89700 582472 89712
rect 582524 89700 582530 89752
rect 582374 86204 582380 86216
rect 582335 86176 582380 86204
rect 582374 86164 582380 86176
rect 582432 86164 582438 86216
rect 582374 75936 582380 75948
rect 582335 75908 582380 75936
rect 582374 75896 582380 75908
rect 582432 75896 582438 75948
rect 582558 73012 582564 73024
rect 582519 72984 582564 73012
rect 582558 72972 582564 72984
rect 582616 72972 582622 73024
rect 582558 60772 582564 60784
rect 582519 60744 582564 60772
rect 582558 60732 582564 60744
rect 582616 60732 582622 60784
rect 582466 59684 582472 59696
rect 582427 59656 582472 59684
rect 582466 59644 582472 59656
rect 582524 59644 582530 59696
rect 582374 46356 582380 46368
rect 582335 46328 582380 46356
rect 582374 46316 582380 46328
rect 582432 46316 582438 46368
rect 582650 46152 582656 46164
rect 582611 46124 582656 46152
rect 582650 46112 582656 46124
rect 582708 46112 582714 46164
rect 582558 33096 582564 33108
rect 582519 33068 582564 33096
rect 582558 33056 582564 33068
rect 582616 33056 582622 33108
rect 582466 31804 582472 31816
rect 582427 31776 582472 31804
rect 582466 31764 582472 31776
rect 582524 31764 582530 31816
rect 303614 29792 303620 29844
rect 303672 29832 303678 29844
rect 304762 29832 304768 29844
rect 303672 29804 304768 29832
rect 303672 29792 303678 29804
rect 304762 29792 304768 29804
rect 304820 29792 304826 29844
rect 318794 29792 318800 29844
rect 318852 29832 318858 29844
rect 319942 29832 319948 29844
rect 318852 29804 319948 29832
rect 318852 29792 318858 29804
rect 319942 29792 319948 29804
rect 320000 29792 320006 29844
rect 333974 29792 333980 29844
rect 334032 29832 334038 29844
rect 335122 29832 335128 29844
rect 334032 29804 335128 29832
rect 334032 29792 334038 29804
rect 335122 29792 335128 29804
rect 335180 29792 335186 29844
rect 349154 29792 349160 29844
rect 349212 29832 349218 29844
rect 350302 29832 350308 29844
rect 349212 29804 350308 29832
rect 349212 29792 349218 29804
rect 350302 29792 350308 29804
rect 350360 29792 350366 29844
rect 379514 29792 379520 29844
rect 379572 29832 379578 29844
rect 380662 29832 380668 29844
rect 379572 29804 380668 29832
rect 379572 29792 379578 29804
rect 380662 29792 380668 29804
rect 380720 29792 380726 29844
rect 425054 29792 425060 29844
rect 425112 29832 425118 29844
rect 426202 29832 426208 29844
rect 425112 29804 426208 29832
rect 425112 29792 425118 29804
rect 426202 29792 426208 29804
rect 426260 29792 426266 29844
rect 440234 29792 440240 29844
rect 440292 29832 440298 29844
rect 441474 29832 441480 29844
rect 440292 29804 441480 29832
rect 440292 29792 440298 29804
rect 441474 29792 441480 29804
rect 441532 29792 441538 29844
rect 470594 29792 470600 29844
rect 470652 29832 470658 29844
rect 471834 29832 471840 29844
rect 470652 29804 471840 29832
rect 470652 29792 470658 29804
rect 471834 29792 471840 29804
rect 471892 29792 471898 29844
rect 500954 29792 500960 29844
rect 501012 29832 501018 29844
rect 502194 29832 502200 29844
rect 501012 29804 502200 29832
rect 501012 29792 501018 29804
rect 502194 29792 502200 29804
rect 502252 29792 502258 29844
rect 561674 29792 561680 29844
rect 561732 29832 561738 29844
rect 562914 29832 562920 29844
rect 561732 29804 562920 29832
rect 561732 29792 561738 29804
rect 562914 29792 562920 29804
rect 562972 29792 562978 29844
rect 1302 27548 1308 27600
rect 1360 27588 1366 27600
rect 5994 27588 6000 27600
rect 1360 27560 6000 27588
rect 1360 27548 1366 27560
rect 5994 27548 6000 27560
rect 6052 27548 6058 27600
rect 26326 27548 26332 27600
rect 26384 27588 26390 27600
rect 29638 27588 29644 27600
rect 26384 27560 29644 27588
rect 26384 27548 26390 27560
rect 29638 27548 29644 27560
rect 29696 27548 29702 27600
rect 36446 27548 36452 27600
rect 36504 27588 36510 27600
rect 39298 27588 39304 27600
rect 36504 27560 39304 27588
rect 36504 27548 36510 27560
rect 39298 27548 39304 27560
rect 39356 27548 39362 27600
rect 41506 27548 41512 27600
rect 41564 27588 41570 27600
rect 43438 27588 43444 27600
rect 41564 27560 43444 27588
rect 41564 27548 41570 27560
rect 43438 27548 43444 27560
rect 43496 27548 43502 27600
rect 46566 27548 46572 27600
rect 46624 27588 46630 27600
rect 47578 27588 47584 27600
rect 46624 27560 47584 27588
rect 46624 27548 46630 27560
rect 47578 27548 47584 27560
rect 47636 27548 47642 27600
rect 51626 27548 51632 27600
rect 51684 27588 51690 27600
rect 52362 27588 52368 27600
rect 51684 27560 52368 27588
rect 51684 27548 51690 27560
rect 52362 27548 52368 27560
rect 52420 27548 52426 27600
rect 56686 27548 56692 27600
rect 56744 27588 56750 27600
rect 57882 27588 57888 27600
rect 56744 27560 57888 27588
rect 56744 27548 56750 27560
rect 57882 27548 57888 27560
rect 57940 27548 57946 27600
rect 58618 27548 58624 27600
rect 58676 27588 58682 27600
rect 122374 27588 122380 27600
rect 58676 27560 122380 27588
rect 58676 27548 58682 27560
rect 122374 27548 122380 27560
rect 122432 27548 122438 27600
rect 124858 27548 124864 27600
rect 124916 27588 124922 27600
rect 127434 27588 127440 27600
rect 124916 27560 127440 27588
rect 124916 27548 124922 27560
rect 127434 27548 127440 27560
rect 127492 27548 127498 27600
rect 162118 27548 162124 27600
rect 162176 27588 162182 27600
rect 162946 27588 162952 27600
rect 162176 27560 162952 27588
rect 162176 27548 162182 27560
rect 162946 27548 162952 27560
rect 163004 27548 163010 27600
rect 166258 27548 166264 27600
rect 166316 27588 166322 27600
rect 168006 27588 168012 27600
rect 166316 27560 168012 27588
rect 166316 27548 166322 27560
rect 168006 27548 168012 27560
rect 168064 27548 168070 27600
rect 190454 27548 190460 27600
rect 190512 27588 190518 27600
rect 193306 27588 193312 27600
rect 190512 27560 193312 27588
rect 190512 27548 190518 27560
rect 193306 27548 193312 27560
rect 193364 27548 193370 27600
rect 313918 27548 313924 27600
rect 313976 27588 313982 27600
rect 314838 27588 314844 27600
rect 313976 27560 314844 27588
rect 313976 27548 313982 27560
rect 314838 27548 314844 27560
rect 314896 27548 314902 27600
rect 454678 27548 454684 27600
rect 454736 27588 454742 27600
rect 456610 27588 456616 27600
rect 454736 27560 456616 27588
rect 454736 27548 454742 27560
rect 456610 27548 456616 27560
rect 456668 27548 456674 27600
rect 53098 27480 53104 27532
rect 53156 27520 53162 27532
rect 132494 27520 132500 27532
rect 53156 27492 132500 27520
rect 53156 27480 53162 27492
rect 132494 27480 132500 27492
rect 132552 27480 132558 27532
rect 66806 27412 66812 27464
rect 66864 27452 66870 27464
rect 69658 27452 69664 27464
rect 66864 27424 69664 27452
rect 66864 27412 66870 27424
rect 69658 27412 69664 27424
rect 69716 27412 69722 27464
rect 81986 27412 81992 27464
rect 82044 27452 82050 27464
rect 83458 27452 83464 27464
rect 82044 27424 83464 27452
rect 82044 27412 82050 27424
rect 83458 27412 83464 27424
rect 83516 27412 83522 27464
rect 83553 27455 83611 27461
rect 83553 27421 83565 27455
rect 83599 27452 83611 27455
rect 97074 27452 97080 27464
rect 83599 27424 97080 27452
rect 83599 27421 83611 27424
rect 83553 27415 83611 27421
rect 97074 27412 97080 27424
rect 97132 27412 97138 27464
rect 101398 27412 101404 27464
rect 101456 27452 101462 27464
rect 102134 27452 102140 27464
rect 101456 27424 102140 27452
rect 101456 27412 101462 27424
rect 102134 27412 102140 27424
rect 102192 27412 102198 27464
rect 114462 27412 114468 27464
rect 114520 27452 114526 27464
rect 365438 27452 365444 27464
rect 114520 27424 365444 27452
rect 114520 27412 114526 27424
rect 365438 27412 365444 27424
rect 365496 27412 365502 27464
rect 68278 27344 68284 27396
rect 68336 27384 68342 27396
rect 107194 27384 107200 27396
rect 68336 27356 107200 27384
rect 68336 27344 68342 27356
rect 107194 27344 107200 27356
rect 107252 27344 107258 27396
rect 107562 27344 107568 27396
rect 107620 27384 107626 27396
rect 375558 27384 375564 27396
rect 107620 27356 375564 27384
rect 107620 27344 107626 27356
rect 375558 27344 375564 27356
rect 375616 27344 375622 27396
rect 71866 27276 71872 27328
rect 71924 27316 71930 27328
rect 90358 27316 90364 27328
rect 71924 27288 90364 27316
rect 71924 27276 71930 27288
rect 90358 27276 90364 27288
rect 90416 27276 90422 27328
rect 93762 27276 93768 27328
rect 93820 27316 93826 27328
rect 395798 27316 395804 27328
rect 93820 27288 395804 27316
rect 93820 27276 93826 27288
rect 395798 27276 395804 27288
rect 395856 27276 395862 27328
rect 75178 27208 75184 27260
rect 75236 27248 75242 27260
rect 83553 27251 83611 27257
rect 83553 27248 83565 27251
rect 75236 27220 83565 27248
rect 75236 27208 75242 27220
rect 83553 27217 83565 27220
rect 83599 27217 83611 27251
rect 83553 27211 83611 27217
rect 86770 27208 86776 27260
rect 86828 27248 86834 27260
rect 405918 27248 405924 27260
rect 86828 27220 405924 27248
rect 86828 27208 86834 27220
rect 405918 27208 405924 27220
rect 405976 27208 405982 27260
rect 31386 27140 31392 27192
rect 31444 27180 31450 27192
rect 50338 27180 50344 27192
rect 31444 27152 50344 27180
rect 31444 27140 31450 27152
rect 50338 27140 50344 27152
rect 50396 27140 50402 27192
rect 82722 27140 82728 27192
rect 82780 27180 82786 27192
rect 410978 27180 410984 27192
rect 82780 27152 410984 27180
rect 82780 27140 82786 27152
rect 410978 27140 410984 27152
rect 411036 27140 411042 27192
rect 486418 27140 486424 27192
rect 486476 27180 486482 27192
rect 486476 27152 489914 27180
rect 486476 27140 486482 27152
rect 33778 27072 33784 27124
rect 33836 27112 33842 27124
rect 486970 27112 486976 27124
rect 33836 27084 486976 27112
rect 33836 27072 33842 27084
rect 486970 27072 486976 27084
rect 487028 27072 487034 27124
rect 489886 27112 489914 27152
rect 527450 27112 527456 27124
rect 489886 27084 527456 27112
rect 527450 27072 527456 27084
rect 527508 27072 527514 27124
rect 5442 27004 5448 27056
rect 5500 27044 5506 27056
rect 11054 27044 11060 27056
rect 5500 27016 11060 27044
rect 5500 27004 5506 27016
rect 11054 27004 11060 27016
rect 11112 27004 11118 27056
rect 32398 27004 32404 27056
rect 32456 27044 32462 27056
rect 497090 27044 497096 27056
rect 32456 27016 497096 27044
rect 32456 27004 32462 27016
rect 497090 27004 497096 27016
rect 497148 27004 497154 27056
rect 497458 27004 497464 27056
rect 497516 27044 497522 27056
rect 517330 27044 517336 27056
rect 497516 27016 517336 27044
rect 497516 27004 497522 27016
rect 517330 27004 517336 27016
rect 517388 27004 517394 27056
rect 518158 27004 518164 27056
rect 518216 27044 518222 27056
rect 532510 27044 532516 27056
rect 518216 27016 532516 27044
rect 518216 27004 518222 27016
rect 532510 27004 532516 27016
rect 532568 27004 532574 27056
rect 4062 26936 4068 26988
rect 4120 26976 4126 26988
rect 16114 26976 16120 26988
rect 4120 26948 16120 26976
rect 4120 26936 4126 26948
rect 16114 26936 16120 26948
rect 16172 26936 16178 26988
rect 36538 26936 36544 26988
rect 36596 26976 36602 26988
rect 567930 26976 567936 26988
rect 36596 26948 567936 26976
rect 36596 26936 36602 26948
rect 567930 26936 567936 26948
rect 567988 26936 567994 26988
rect 6822 26868 6828 26920
rect 6880 26908 6886 26920
rect 21174 26908 21180 26920
rect 6880 26880 21180 26908
rect 6880 26868 6886 26880
rect 21174 26868 21180 26880
rect 21232 26868 21238 26920
rect 35158 26868 35164 26920
rect 35216 26908 35222 26920
rect 578142 26908 578148 26920
rect 35216 26880 578148 26908
rect 35216 26868 35222 26880
rect 578142 26868 578148 26880
rect 578200 26868 578206 26920
rect 65518 26800 65524 26852
rect 65576 26840 65582 26852
rect 117314 26840 117320 26852
rect 65576 26812 117320 26840
rect 65576 26800 65582 26812
rect 117314 26800 117320 26812
rect 117372 26800 117378 26852
rect 79318 26732 79324 26784
rect 79376 26772 79382 26784
rect 92014 26772 92020 26784
rect 79376 26744 92020 26772
rect 79376 26732 79382 26744
rect 92014 26732 92020 26744
rect 92072 26732 92078 26784
rect 40678 25712 40684 25764
rect 40736 25752 40742 25764
rect 157334 25752 157340 25764
rect 40736 25724 157340 25752
rect 40736 25712 40742 25724
rect 157334 25712 157340 25724
rect 157392 25712 157398 25764
rect 18598 25644 18604 25696
rect 18656 25684 18662 25696
rect 182174 25684 182180 25696
rect 18656 25656 182180 25684
rect 18656 25644 18662 25656
rect 182174 25644 182180 25656
rect 182232 25644 182238 25696
rect 54478 25576 54484 25628
rect 54536 25616 54542 25628
rect 451274 25616 451280 25628
rect 54536 25588 451280 25616
rect 54536 25576 54542 25588
rect 451274 25576 451280 25588
rect 451332 25576 451338 25628
rect 7558 25508 7564 25560
rect 7616 25548 7622 25560
rect 552014 25548 552020 25560
rect 7616 25520 552020 25548
rect 7616 25508 7622 25520
rect 552014 25508 552020 25520
rect 552072 25508 552078 25560
rect 11698 24080 11704 24132
rect 11756 24120 11762 24132
rect 506474 24120 506480 24132
rect 11756 24092 506480 24120
rect 11756 24080 11762 24092
rect 506474 24080 506480 24092
rect 506532 24080 506538 24132
rect 119982 22720 119988 22772
rect 120040 22760 120046 22772
rect 190454 22760 190460 22772
rect 120040 22732 190460 22760
rect 120040 22720 120046 22732
rect 190454 22720 190460 22732
rect 190512 22720 190518 22772
rect 29638 21360 29644 21412
rect 29696 21400 29702 21412
rect 122834 21400 122840 21412
rect 29696 21372 122840 21400
rect 29696 21360 29702 21372
rect 122834 21360 122840 21372
rect 122892 21360 122898 21412
rect 25498 19932 25504 19984
rect 25556 19972 25562 19984
rect 172514 19972 172520 19984
rect 25556 19944 172520 19972
rect 25556 19932 25562 19944
rect 172514 19932 172520 19944
rect 172572 19932 172578 19984
rect 582650 19836 582656 19848
rect 582611 19808 582656 19836
rect 582650 19796 582656 19808
rect 582708 19796 582714 19848
rect 62022 18572 62028 18624
rect 62080 18612 62086 18624
rect 97994 18612 98000 18624
rect 62080 18584 98000 18612
rect 62080 18572 62086 18584
rect 97994 18572 98000 18584
rect 98052 18572 98058 18624
rect 52362 17212 52368 17264
rect 52420 17252 52426 17264
rect 104894 17252 104900 17264
rect 52420 17224 104900 17252
rect 52420 17212 52426 17224
rect 104894 17212 104900 17224
rect 104952 17212 104958 17264
rect 69658 15920 69664 15972
rect 69716 15960 69722 15972
rect 94682 15960 94688 15972
rect 69716 15932 94688 15960
rect 69716 15920 69722 15932
rect 94682 15920 94688 15932
rect 94740 15920 94746 15972
rect 51718 15852 51724 15904
rect 51776 15892 51782 15904
rect 142154 15892 142160 15904
rect 51776 15864 142160 15892
rect 51776 15852 51782 15864
rect 142154 15852 142160 15864
rect 142212 15852 142218 15904
rect 144730 15852 144736 15904
rect 144788 15892 144794 15904
rect 536834 15892 536840 15904
rect 144788 15864 536840 15892
rect 144788 15852 144794 15864
rect 536834 15852 536840 15864
rect 536892 15852 536898 15904
rect 41322 14424 41328 14476
rect 41380 14464 41386 14476
rect 303614 14464 303620 14476
rect 41380 14436 303620 14464
rect 41380 14424 41386 14436
rect 303614 14424 303620 14436
rect 303672 14424 303678 14476
rect 22738 13064 22744 13116
rect 22796 13104 22802 13116
rect 178034 13104 178040 13116
rect 22796 13076 178040 13104
rect 22796 13064 22802 13076
rect 178034 13064 178040 13076
rect 178092 13064 178098 13116
rect 70302 11772 70308 11824
rect 70360 11812 70366 11824
rect 101398 11812 101404 11824
rect 70360 11784 101404 11812
rect 70360 11772 70366 11784
rect 101398 11772 101404 11784
rect 101456 11772 101462 11824
rect 39298 11704 39304 11756
rect 39356 11744 39362 11756
rect 116394 11744 116400 11756
rect 39356 11716 116400 11744
rect 39356 11704 39362 11716
rect 116394 11704 116400 11716
rect 116452 11704 116458 11756
rect 125870 11704 125876 11756
rect 125928 11744 125934 11756
rect 486418 11744 486424 11756
rect 125928 11716 486424 11744
rect 125928 11704 125934 11716
rect 486418 11704 486424 11716
rect 486476 11704 486482 11756
rect 39298 10344 39304 10396
rect 39356 10384 39362 10396
rect 151814 10384 151820 10396
rect 39356 10356 151820 10384
rect 39356 10344 39362 10356
rect 151814 10344 151820 10356
rect 151872 10344 151878 10396
rect 14458 10276 14464 10328
rect 14516 10316 14522 10328
rect 557534 10316 557540 10328
rect 14516 10288 557540 10316
rect 14516 10276 14522 10288
rect 557534 10276 557540 10288
rect 557592 10276 557598 10328
rect 27706 9120 27712 9172
rect 27764 9160 27770 9172
rect 162118 9160 162124 9172
rect 27764 9132 162124 9160
rect 27764 9120 27770 9132
rect 162118 9120 162124 9132
rect 162176 9120 162182 9172
rect 44266 9052 44272 9104
rect 44324 9092 44330 9104
rect 299474 9092 299480 9104
rect 44324 9064 299480 9092
rect 44324 9052 44330 9064
rect 299474 9052 299480 9064
rect 299532 9052 299538 9104
rect 49878 8984 49884 9036
rect 49936 9024 49942 9036
rect 136634 9024 136640 9036
rect 49936 8996 136640 9024
rect 49936 8984 49942 8996
rect 136634 8984 136640 8996
rect 136692 8984 136698 9036
rect 141234 8984 141240 9036
rect 141292 9024 141298 9036
rect 542354 9024 542360 9036
rect 141292 8996 542360 9024
rect 141292 8984 141298 8996
rect 542354 8984 542360 8996
rect 542412 8984 542418 9036
rect 50154 8916 50160 8968
rect 50212 8956 50218 8968
rect 454678 8956 454684 8968
rect 50212 8928 454684 8956
rect 50212 8916 50218 8928
rect 454678 8916 454684 8928
rect 454736 8916 454742 8968
rect 122282 7964 122288 8016
rect 122340 8004 122346 8016
rect 187694 8004 187700 8016
rect 122340 7976 187700 8004
rect 122340 7964 122346 7976
rect 187694 7964 187700 7976
rect 187752 7964 187758 8016
rect 23014 7896 23020 7948
rect 23072 7936 23078 7948
rect 166258 7936 166264 7948
rect 23072 7908 166264 7936
rect 23072 7896 23078 7908
rect 166258 7896 166264 7908
rect 166316 7896 166322 7948
rect 37182 7828 37188 7880
rect 37240 7868 37246 7880
rect 309134 7868 309140 7880
rect 37240 7840 309140 7868
rect 37240 7828 37246 7840
rect 309134 7828 309140 7840
rect 309192 7828 309198 7880
rect 33594 7760 33600 7812
rect 33652 7800 33658 7812
rect 313918 7800 313924 7812
rect 33652 7772 313924 7800
rect 33652 7760 33658 7772
rect 313918 7760 313924 7772
rect 313976 7760 313982 7812
rect 50338 7692 50344 7744
rect 50396 7732 50402 7744
rect 119890 7732 119896 7744
rect 50396 7704 119896 7732
rect 50396 7692 50402 7704
rect 119890 7692 119896 7704
rect 119948 7692 119954 7744
rect 132954 7692 132960 7744
rect 133012 7732 133018 7744
rect 497458 7732 497464 7744
rect 133012 7704 497464 7732
rect 133012 7692 133018 7704
rect 497458 7692 497464 7704
rect 497516 7692 497522 7744
rect 43162 7624 43168 7676
rect 43220 7664 43226 7676
rect 147674 7664 147680 7676
rect 43220 7636 147680 7664
rect 43220 7624 43226 7636
rect 147674 7624 147680 7636
rect 147732 7624 147738 7676
rect 148318 7624 148324 7676
rect 148376 7664 148382 7676
rect 518158 7664 518164 7676
rect 148376 7636 518164 7664
rect 148376 7624 148382 7636
rect 518158 7624 518164 7636
rect 518216 7624 518222 7676
rect 43438 7556 43444 7608
rect 43496 7596 43502 7608
rect 112806 7596 112812 7608
rect 43496 7568 112812 7596
rect 43496 7556 43502 7568
rect 112806 7556 112812 7568
rect 112864 7556 112870 7608
rect 129366 7556 129372 7608
rect 129424 7596 129430 7608
rect 521654 7596 521660 7608
rect 129424 7568 521660 7596
rect 129424 7556 129430 7568
rect 521654 7556 521660 7568
rect 521712 7556 521718 7608
rect 80882 6808 80888 6860
rect 80940 6848 80946 6860
rect 86954 6848 86960 6860
rect 80940 6820 86960 6848
rect 80940 6808 80946 6820
rect 86954 6808 86960 6820
rect 87012 6808 87018 6860
rect 77202 6672 77208 6724
rect 77260 6712 77266 6724
rect 87966 6712 87972 6724
rect 77260 6684 87972 6712
rect 77260 6672 77266 6684
rect 87966 6672 87972 6684
rect 88024 6672 88030 6724
rect 63218 6604 63224 6656
rect 63276 6644 63282 6656
rect 111794 6644 111800 6656
rect 63276 6616 111800 6644
rect 63276 6604 63282 6616
rect 111794 6604 111800 6616
rect 111852 6604 111858 6656
rect 115198 6604 115204 6656
rect 115256 6644 115262 6656
rect 197354 6644 197360 6656
rect 115256 6616 197360 6644
rect 115256 6604 115262 6616
rect 197354 6604 197360 6616
rect 197412 6604 197418 6656
rect 582466 6644 582472 6656
rect 582427 6616 582472 6644
rect 582466 6604 582472 6616
rect 582524 6604 582530 6656
rect 47578 6536 47584 6588
rect 47636 6576 47642 6588
rect 109310 6576 109316 6588
rect 47636 6548 109316 6576
rect 47636 6536 47642 6548
rect 109310 6536 109316 6548
rect 109368 6536 109374 6588
rect 111610 6536 111616 6588
rect 111668 6576 111674 6588
rect 202874 6576 202880 6588
rect 111668 6548 202880 6576
rect 111668 6536 111674 6548
rect 202874 6536 202880 6548
rect 202932 6536 202938 6588
rect 57882 6468 57888 6520
rect 57940 6508 57946 6520
rect 102226 6508 102232 6520
rect 57940 6480 102232 6508
rect 57940 6468 57946 6480
rect 102226 6468 102232 6480
rect 102284 6468 102290 6520
rect 108114 6468 108120 6520
rect 108172 6508 108178 6520
rect 208394 6508 208400 6520
rect 108172 6480 208400 6508
rect 108172 6468 108178 6480
rect 208394 6468 208400 6480
rect 208452 6468 208458 6520
rect 30098 6400 30104 6452
rect 30156 6440 30162 6452
rect 318794 6440 318800 6452
rect 30156 6412 318800 6440
rect 30156 6400 30162 6412
rect 318794 6400 318800 6412
rect 318852 6400 318858 6452
rect 26510 6332 26516 6384
rect 26568 6372 26574 6384
rect 324314 6372 324320 6384
rect 26568 6344 324320 6372
rect 26568 6332 26574 6344
rect 324314 6332 324320 6344
rect 324372 6332 324378 6384
rect 21818 6264 21824 6316
rect 21876 6304 21882 6316
rect 329834 6304 329840 6316
rect 21876 6276 329840 6304
rect 21876 6264 21882 6276
rect 329834 6264 329840 6276
rect 329892 6264 329898 6316
rect 17034 6196 17040 6248
rect 17092 6236 17098 6248
rect 333974 6236 333980 6248
rect 17092 6208 333980 6236
rect 17092 6196 17098 6208
rect 333974 6196 333980 6208
rect 334032 6196 334038 6248
rect 52546 6128 52552 6180
rect 52604 6168 52610 6180
rect 124858 6168 124864 6180
rect 52604 6140 124864 6168
rect 52604 6128 52610 6140
rect 124858 6128 124864 6140
rect 124916 6128 124922 6180
rect 136450 6128 136456 6180
rect 136508 6168 136514 6180
rect 511994 6168 512000 6180
rect 136508 6140 512000 6168
rect 136508 6128 136514 6140
rect 511994 6128 512000 6140
rect 512052 6128 512058 6180
rect 76190 5448 76196 5500
rect 76248 5488 76254 5500
rect 253934 5488 253940 5500
rect 76248 5460 253940 5488
rect 76248 5448 76254 5460
rect 253934 5448 253940 5460
rect 253992 5448 253998 5500
rect 72602 5380 72608 5432
rect 72660 5420 72666 5432
rect 258074 5420 258080 5432
rect 72660 5392 258080 5420
rect 72660 5380 72666 5392
rect 258074 5380 258080 5392
rect 258132 5380 258138 5432
rect 69106 5312 69112 5364
rect 69164 5352 69170 5364
rect 263594 5352 263600 5364
rect 69164 5324 263600 5352
rect 69164 5312 69170 5324
rect 263594 5312 263600 5324
rect 263652 5312 263658 5364
rect 65610 5244 65616 5296
rect 65668 5284 65674 5296
rect 269114 5284 269120 5296
rect 65668 5256 269120 5284
rect 65668 5244 65674 5256
rect 269114 5244 269120 5256
rect 269172 5244 269178 5296
rect 62022 5176 62028 5228
rect 62080 5216 62086 5228
rect 273254 5216 273260 5228
rect 62080 5188 273260 5216
rect 62080 5176 62086 5188
rect 273254 5176 273260 5188
rect 273312 5176 273318 5228
rect 58434 5108 58440 5160
rect 58492 5148 58498 5160
rect 278774 5148 278780 5160
rect 58492 5120 278780 5148
rect 58492 5108 58498 5120
rect 278774 5108 278780 5120
rect 278832 5108 278838 5160
rect 54938 5040 54944 5092
rect 54996 5080 55002 5092
rect 284294 5080 284300 5092
rect 54996 5052 284300 5080
rect 54996 5040 55002 5052
rect 284294 5040 284300 5052
rect 284352 5040 284358 5092
rect 51350 4972 51356 5024
rect 51408 5012 51414 5024
rect 288434 5012 288440 5024
rect 51408 4984 288440 5012
rect 51408 4972 51414 4984
rect 288434 4972 288440 4984
rect 288492 4972 288498 5024
rect 47854 4904 47860 4956
rect 47912 4944 47918 4956
rect 293954 4944 293960 4956
rect 47912 4916 293960 4944
rect 47912 4904 47918 4916
rect 293954 4904 293960 4916
rect 294012 4904 294018 4956
rect 12342 4836 12348 4888
rect 12400 4876 12406 4888
rect 339494 4876 339500 4888
rect 12400 4848 339500 4876
rect 12400 4836 12406 4848
rect 339494 4836 339500 4848
rect 339552 4836 339558 4888
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 345014 4808 345020 4820
rect 7708 4780 345020 4808
rect 7708 4768 7714 4780
rect 345014 4768 345020 4780
rect 345072 4768 345078 4820
rect 73798 4700 73804 4752
rect 73856 4740 73862 4752
rect 75178 4740 75184 4752
rect 73856 4712 75184 4740
rect 73856 4700 73862 4712
rect 75178 4700 75184 4712
rect 75236 4700 75242 4752
rect 83458 4700 83464 4752
rect 83516 4740 83522 4752
rect 84470 4740 84476 4752
rect 83516 4712 84476 4740
rect 83516 4700 83522 4712
rect 84470 4700 84476 4712
rect 84528 4700 84534 4752
rect 248414 4740 248420 4752
rect 88996 4712 248420 4740
rect 79686 4564 79692 4616
rect 79744 4604 79750 4616
rect 88996 4604 89024 4712
rect 248414 4700 248420 4712
rect 248472 4700 248478 4752
rect 242894 4672 242900 4684
rect 79744 4576 89024 4604
rect 89088 4644 242900 4672
rect 79744 4564 79750 4576
rect 83274 4496 83280 4548
rect 83332 4536 83338 4548
rect 89088 4536 89116 4644
rect 242894 4632 242900 4644
rect 242952 4632 242958 4684
rect 238754 4604 238760 4616
rect 83332 4508 89116 4536
rect 89180 4576 238760 4604
rect 83332 4496 83338 4508
rect 86862 4428 86868 4480
rect 86920 4468 86926 4480
rect 89180 4468 89208 4576
rect 238754 4564 238760 4576
rect 238812 4564 238818 4616
rect 90450 4496 90456 4548
rect 90508 4536 90514 4548
rect 233234 4536 233240 4548
rect 90508 4508 233240 4536
rect 90508 4496 90514 4508
rect 233234 4496 233240 4508
rect 233292 4496 233298 4548
rect 86920 4440 89208 4468
rect 86920 4428 86926 4440
rect 93946 4428 93952 4480
rect 94004 4468 94010 4480
rect 227714 4468 227720 4480
rect 94004 4440 227720 4468
rect 94004 4428 94010 4440
rect 227714 4428 227720 4440
rect 227772 4428 227778 4480
rect 59630 4360 59636 4412
rect 59688 4400 59694 4412
rect 65518 4400 65524 4412
rect 59688 4372 65524 4400
rect 59688 4360 59694 4372
rect 65518 4360 65524 4372
rect 65576 4360 65582 4412
rect 97442 4360 97448 4412
rect 97500 4400 97506 4412
rect 223574 4400 223580 4412
rect 97500 4372 223580 4400
rect 97500 4360 97506 4372
rect 223574 4360 223580 4372
rect 223632 4360 223638 4412
rect 101030 4292 101036 4344
rect 101088 4332 101094 4344
rect 218054 4332 218060 4344
rect 101088 4304 218060 4332
rect 101088 4292 101094 4304
rect 218054 4292 218060 4304
rect 218112 4292 218118 4344
rect 104526 4224 104532 4276
rect 104584 4264 104590 4276
rect 212534 4264 212540 4276
rect 104584 4236 212540 4264
rect 104584 4224 104590 4236
rect 212534 4224 212540 4236
rect 212592 4224 212598 4276
rect 48958 4156 48964 4208
rect 49016 4196 49022 4208
rect 53098 4196 53104 4208
rect 49016 4168 53104 4196
rect 49016 4156 49022 4168
rect 53098 4156 53104 4168
rect 53156 4156 53162 4208
rect 56042 4156 56048 4208
rect 56100 4196 56106 4208
rect 58618 4196 58624 4208
rect 56100 4168 58624 4196
rect 56100 4156 56106 4168
rect 58618 4156 58624 4168
rect 58676 4156 58682 4208
rect 66714 4156 66720 4208
rect 66772 4196 66778 4208
rect 68278 4196 68284 4208
rect 66772 4168 68284 4196
rect 66772 4156 66778 4168
rect 68278 4156 68284 4168
rect 68336 4156 68342 4208
rect 77386 4156 77392 4208
rect 77444 4196 77450 4208
rect 79318 4196 79324 4208
rect 77444 4168 79324 4196
rect 77444 4156 77450 4168
rect 79318 4156 79324 4168
rect 79376 4156 79382 4208
rect 90358 4156 90364 4208
rect 90416 4196 90422 4208
rect 91554 4196 91560 4208
rect 90416 4168 91560 4196
rect 90416 4156 90422 4168
rect 91554 4156 91560 4168
rect 91612 4156 91618 4208
rect 1670 4088 1676 4140
rect 1728 4128 1734 4140
rect 7558 4128 7564 4140
rect 1728 4100 7564 4128
rect 1728 4088 1734 4100
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 74994 4088 75000 4140
rect 75052 4128 75058 4140
rect 420914 4128 420920 4140
rect 75052 4100 420920 4128
rect 75052 4088 75058 4100
rect 420914 4088 420920 4100
rect 420972 4088 420978 4140
rect 71498 4020 71504 4072
rect 71556 4060 71562 4072
rect 425054 4060 425060 4072
rect 71556 4032 425060 4060
rect 71556 4020 71562 4032
rect 425054 4020 425060 4032
rect 425112 4020 425118 4072
rect 67910 3952 67916 4004
rect 67968 3992 67974 4004
rect 430574 3992 430580 4004
rect 67968 3964 430580 3992
rect 67968 3952 67974 3964
rect 430574 3952 430580 3964
rect 430632 3952 430638 4004
rect 64322 3884 64328 3936
rect 64380 3924 64386 3936
rect 436094 3924 436100 3936
rect 64380 3896 436100 3924
rect 64380 3884 64386 3896
rect 436094 3884 436100 3896
rect 436152 3884 436158 3936
rect 45462 3816 45468 3868
rect 45520 3856 45526 3868
rect 49878 3856 49884 3868
rect 45520 3828 49884 3856
rect 45520 3816 45526 3828
rect 49878 3816 49884 3828
rect 49936 3816 49942 3868
rect 60826 3816 60832 3868
rect 60884 3856 60890 3868
rect 440234 3856 440240 3868
rect 60884 3828 440240 3856
rect 60884 3816 60890 3828
rect 440234 3816 440240 3828
rect 440292 3816 440298 3868
rect 41874 3748 41880 3800
rect 41932 3788 41938 3800
rect 51718 3788 51724 3800
rect 41932 3760 51724 3788
rect 41932 3748 41938 3760
rect 51718 3748 51724 3760
rect 51776 3748 51782 3800
rect 57238 3748 57244 3800
rect 57296 3788 57302 3800
rect 445754 3788 445760 3800
rect 57296 3760 445760 3788
rect 57296 3748 57302 3760
rect 445754 3748 445760 3760
rect 445812 3748 445818 3800
rect 13538 3680 13544 3732
rect 13596 3720 13602 3732
rect 22738 3720 22744 3732
rect 13596 3692 22744 3720
rect 13596 3680 13602 3692
rect 22738 3680 22744 3692
rect 22796 3680 22802 3732
rect 31294 3680 31300 3732
rect 31352 3720 31358 3732
rect 40678 3720 40684 3732
rect 31352 3692 40684 3720
rect 31352 3680 31358 3692
rect 40678 3680 40684 3692
rect 40736 3680 40742 3732
rect 46658 3680 46664 3732
rect 46716 3720 46722 3732
rect 460934 3720 460940 3732
rect 46716 3692 460940 3720
rect 46716 3680 46722 3692
rect 460934 3680 460940 3692
rect 460992 3680 460998 3732
rect 19426 3612 19432 3664
rect 19484 3652 19490 3664
rect 32398 3652 32404 3664
rect 19484 3624 32404 3652
rect 19484 3612 19490 3624
rect 32398 3612 32404 3624
rect 32456 3612 32462 3664
rect 34790 3612 34796 3664
rect 34848 3652 34854 3664
rect 39298 3652 39304 3664
rect 34848 3624 39304 3652
rect 34848 3612 34854 3624
rect 39298 3612 39304 3624
rect 39356 3612 39362 3664
rect 43070 3612 43076 3664
rect 43128 3652 43134 3664
rect 466454 3652 466460 3664
rect 43128 3624 466460 3652
rect 43128 3612 43134 3624
rect 466454 3612 466460 3624
rect 466512 3612 466518 3664
rect 8754 3544 8760 3596
rect 8812 3584 8818 3596
rect 18598 3584 18604 3596
rect 8812 3556 18604 3584
rect 8812 3544 8818 3556
rect 18598 3544 18604 3556
rect 18656 3544 18662 3596
rect 20622 3544 20628 3596
rect 20680 3584 20686 3596
rect 36538 3584 36544 3596
rect 20680 3556 36544 3584
rect 20680 3544 20686 3556
rect 36538 3544 36544 3556
rect 36596 3544 36602 3596
rect 39574 3544 39580 3596
rect 39632 3584 39638 3596
rect 470594 3584 470600 3596
rect 39632 3556 470600 3584
rect 39632 3544 39638 3556
rect 470594 3544 470600 3556
rect 470652 3544 470658 3596
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 1302 3516 1308 3528
rect 624 3488 1308 3516
rect 624 3476 630 3488
rect 1302 3476 1308 3488
rect 1360 3476 1366 3528
rect 11146 3476 11152 3528
rect 11204 3516 11210 3528
rect 11204 3488 26234 3516
rect 11204 3476 11210 3488
rect 2866 3408 2872 3460
rect 2924 3448 2930 3460
rect 14458 3448 14464 3460
rect 2924 3420 14464 3448
rect 2924 3408 2930 3420
rect 14458 3408 14464 3420
rect 14516 3408 14522 3460
rect 26206 3448 26234 3488
rect 28902 3476 28908 3528
rect 28960 3516 28966 3528
rect 33778 3516 33784 3528
rect 28960 3488 33784 3516
rect 28960 3476 28966 3488
rect 33778 3476 33784 3488
rect 33836 3476 33842 3528
rect 40678 3476 40684 3528
rect 40736 3516 40742 3528
rect 41322 3516 41328 3528
rect 40736 3488 41328 3516
rect 40736 3476 40742 3488
rect 41322 3476 41328 3488
rect 41380 3476 41386 3528
rect 476114 3516 476120 3528
rect 41524 3488 476120 3516
rect 35158 3448 35164 3460
rect 26206 3420 35164 3448
rect 35158 3408 35164 3420
rect 35216 3408 35222 3460
rect 35986 3340 35992 3392
rect 36044 3380 36050 3392
rect 41524 3380 41552 3488
rect 476114 3476 476120 3488
rect 476172 3476 476178 3528
rect 53742 3408 53748 3460
rect 53800 3448 53806 3460
rect 54478 3448 54484 3460
rect 53800 3420 54484 3448
rect 53800 3408 53806 3420
rect 54478 3408 54484 3420
rect 54536 3408 54542 3460
rect 481634 3448 481640 3460
rect 55186 3420 481640 3448
rect 36044 3352 41552 3380
rect 36044 3340 36050 3352
rect 38378 3272 38384 3324
rect 38436 3312 38442 3324
rect 43162 3312 43168 3324
rect 38436 3284 43168 3312
rect 38436 3272 38442 3284
rect 43162 3272 43168 3284
rect 43220 3272 43226 3324
rect 32398 3204 32404 3256
rect 32456 3244 32462 3256
rect 55186 3244 55214 3420
rect 481634 3408 481640 3420
rect 481692 3408 481698 3460
rect 547782 3408 547788 3460
rect 547840 3448 547846 3460
rect 579798 3448 579804 3460
rect 547840 3420 579804 3448
rect 547840 3408 547846 3420
rect 579798 3408 579804 3420
rect 579856 3408 579862 3460
rect 82078 3340 82084 3392
rect 82136 3380 82142 3392
rect 82722 3380 82728 3392
rect 82136 3352 82728 3380
rect 82136 3340 82142 3352
rect 82722 3340 82728 3352
rect 82780 3340 82786 3392
rect 85666 3340 85672 3392
rect 85724 3380 85730 3392
rect 86770 3380 86776 3392
rect 85724 3352 86776 3380
rect 85724 3340 85730 3352
rect 86770 3340 86776 3352
rect 86828 3340 86834 3392
rect 415394 3380 415400 3392
rect 88996 3352 415400 3380
rect 78582 3272 78588 3324
rect 78640 3312 78646 3324
rect 88996 3312 89024 3352
rect 415394 3340 415400 3352
rect 415452 3340 415458 3392
rect 78640 3284 89024 3312
rect 78640 3272 78646 3284
rect 92750 3272 92756 3324
rect 92808 3312 92814 3324
rect 93762 3312 93768 3324
rect 92808 3284 93768 3312
rect 92808 3272 92814 3284
rect 93762 3272 93768 3284
rect 93820 3272 93826 3324
rect 400214 3312 400220 3324
rect 97828 3284 400220 3312
rect 32456 3216 55214 3244
rect 32456 3204 32462 3216
rect 89162 3204 89168 3256
rect 89220 3244 89226 3256
rect 97828 3244 97856 3284
rect 400214 3272 400220 3284
rect 400272 3272 400278 3324
rect 390554 3244 390560 3256
rect 89220 3216 97856 3244
rect 97920 3216 390560 3244
rect 89220 3204 89226 3216
rect 96246 3136 96252 3188
rect 96304 3176 96310 3188
rect 97920 3176 97948 3216
rect 390554 3204 390560 3216
rect 390612 3204 390618 3256
rect 96304 3148 97948 3176
rect 96304 3136 96310 3148
rect 99834 3136 99840 3188
rect 99892 3176 99898 3188
rect 385034 3176 385040 3188
rect 99892 3148 385040 3176
rect 99892 3136 99898 3148
rect 385034 3136 385040 3148
rect 385092 3136 385098 3188
rect 18230 3068 18236 3120
rect 18288 3108 18294 3120
rect 25498 3108 25504 3120
rect 18288 3080 25504 3108
rect 18288 3068 18294 3080
rect 25498 3068 25504 3080
rect 25556 3068 25562 3120
rect 103330 3068 103336 3120
rect 103388 3108 103394 3120
rect 379514 3108 379520 3120
rect 103388 3080 379520 3108
rect 103388 3068 103394 3080
rect 379514 3068 379520 3080
rect 379572 3068 379578 3120
rect 106918 3000 106924 3052
rect 106976 3040 106982 3052
rect 107562 3040 107568 3052
rect 106976 3012 107568 3040
rect 106976 3000 106982 3012
rect 107562 3000 107568 3012
rect 107620 3000 107626 3052
rect 110506 3000 110512 3052
rect 110564 3040 110570 3052
rect 369854 3040 369860 3052
rect 110564 3012 369860 3040
rect 110564 3000 110570 3012
rect 369854 3000 369860 3012
rect 369912 3000 369918 3052
rect 9950 2932 9956 2984
rect 10008 2972 10014 2984
rect 11698 2972 11704 2984
rect 10008 2944 11704 2972
rect 10008 2932 10014 2944
rect 11698 2932 11704 2944
rect 11756 2932 11762 2984
rect 114002 2932 114008 2984
rect 114060 2972 114066 2984
rect 114462 2972 114468 2984
rect 114060 2944 114468 2972
rect 114060 2932 114066 2944
rect 114462 2932 114468 2944
rect 114520 2932 114526 2984
rect 118786 2932 118792 2984
rect 118844 2972 118850 2984
rect 119982 2972 119988 2984
rect 118844 2944 119988 2972
rect 118844 2932 118850 2944
rect 119982 2932 119988 2944
rect 120040 2932 120046 2984
rect 360194 2972 360200 2984
rect 120092 2944 360200 2972
rect 117590 2864 117596 2916
rect 117648 2904 117654 2916
rect 120092 2904 120120 2944
rect 360194 2932 360200 2944
rect 360252 2932 360258 2984
rect 117648 2876 120120 2904
rect 117648 2864 117654 2876
rect 121086 2864 121092 2916
rect 121144 2904 121150 2916
rect 354674 2904 354680 2916
rect 121144 2876 354680 2904
rect 121144 2864 121150 2876
rect 354674 2864 354680 2876
rect 354732 2864 354738 2916
rect 124674 2796 124680 2848
rect 124732 2836 124738 2848
rect 349154 2836 349160 2848
rect 124732 2808 349160 2836
rect 124732 2796 124738 2808
rect 349154 2796 349160 2808
rect 349212 2796 349218 2848
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 364984 700476 365036 700528
rect 365628 700476 365680 700528
rect 527180 700476 527232 700528
rect 528468 700476 528520 700528
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 105452 700340 105504 700392
rect 106188 700340 106240 700392
rect 235172 700340 235224 700392
rect 235908 700340 235960 700392
rect 170312 700204 170364 700256
rect 171048 700204 171100 700256
rect 397460 699932 397512 699984
rect 398748 699932 398800 699984
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 300124 699660 300176 699712
rect 300768 699660 300820 699712
rect 429844 699660 429896 699712
rect 430488 699660 430540 699712
rect 462320 699660 462372 699712
rect 463608 699660 463660 699712
rect 494796 699660 494848 699712
rect 495348 699660 495400 699712
rect 559656 699660 559708 699712
rect 560208 699660 560260 699712
rect 582380 697187 582432 697196
rect 582380 697153 582389 697187
rect 582389 697153 582423 697187
rect 582423 697153 582432 697187
rect 582380 697144 582432 697153
rect 582472 683859 582524 683868
rect 582472 683825 582481 683859
rect 582481 683825 582515 683859
rect 582515 683825 582524 683859
rect 582472 683816 582524 683825
rect 6092 681640 6144 681692
rect 6920 681640 6972 681692
rect 24768 681640 24820 681692
rect 27988 681640 28040 681692
rect 89628 681640 89680 681692
rect 93952 681640 94004 681692
rect 267648 681232 267700 681284
rect 270040 681232 270092 681284
rect 332508 681096 332560 681148
rect 336004 681096 336056 681148
rect 41328 680960 41380 681012
rect 49976 680960 50028 681012
rect 106188 680960 106240 681012
rect 115940 680960 115992 681012
rect 171048 680960 171100 681012
rect 181996 680960 182048 681012
rect 219348 680960 219400 681012
rect 225972 680960 226024 681012
rect 235908 680960 235960 681012
rect 248052 680960 248104 681012
rect 284208 680960 284260 681012
rect 292028 680960 292080 681012
rect 300768 680960 300820 681012
rect 314016 680960 314068 681012
rect 349068 680960 349120 681012
rect 358084 680960 358136 681012
rect 365628 680960 365680 681012
rect 380072 680960 380124 681012
rect 413928 680960 413980 681012
rect 424048 680960 424100 681012
rect 430488 680960 430540 681012
rect 446036 680960 446088 681012
rect 478788 680960 478840 681012
rect 490104 680960 490156 681012
rect 495348 680960 495400 681012
rect 512092 680960 512144 681012
rect 528468 680960 528520 681012
rect 534080 680960 534132 681012
rect 543648 680960 543700 681012
rect 556068 680960 556120 681012
rect 560208 680960 560260 681012
rect 578056 680960 578108 681012
rect 202788 680892 202840 680944
rect 203984 680892 204036 680944
rect 463608 680892 463660 680944
rect 468116 680892 468168 680944
rect 398748 680688 398800 680740
rect 402060 680688 402112 680740
rect 154488 680620 154540 680672
rect 160008 680620 160060 680672
rect 582380 677535 582432 677544
rect 582380 677501 582389 677535
rect 582389 677501 582423 677535
rect 582423 677501 582432 677535
rect 582380 677492 582432 677501
rect 582380 670735 582432 670744
rect 582380 670701 582389 670735
rect 582389 670701 582423 670735
rect 582423 670701 582432 670735
rect 582380 670692 582432 670701
rect 582472 662371 582524 662380
rect 582472 662337 582481 662371
rect 582481 662337 582515 662371
rect 582515 662337 582524 662371
rect 582472 662328 582524 662337
rect 112 658180 164 658232
rect 572 658180 624 658232
rect 582380 648567 582432 648576
rect 582380 648533 582389 648567
rect 582389 648533 582423 648567
rect 582423 648533 582432 648567
rect 582380 648524 582432 648533
rect 582380 644011 582432 644020
rect 582380 643977 582389 644011
rect 582389 643977 582423 644011
rect 582423 643977 582432 644011
rect 582380 643968 582432 643977
rect 582380 633403 582432 633412
rect 582380 633369 582389 633403
rect 582389 633369 582423 633403
rect 582423 633369 582432 633403
rect 582380 633360 582432 633369
rect 20 632068 72 632120
rect 572 632068 624 632120
rect 582380 630819 582432 630828
rect 582380 630785 582389 630819
rect 582389 630785 582423 630819
rect 582423 630785 582432 630819
rect 582380 630776 582432 630785
rect 582380 618239 582432 618248
rect 582380 618205 582389 618239
rect 582389 618205 582423 618239
rect 582423 618205 582432 618239
rect 582380 618196 582432 618205
rect 582380 617491 582432 617500
rect 582380 617457 582389 617491
rect 582389 617457 582423 617491
rect 582423 617457 582432 617491
rect 582380 617448 582432 617457
rect 582380 604435 582432 604444
rect 582380 604401 582389 604435
rect 582389 604401 582423 604435
rect 582423 604401 582432 604435
rect 582380 604392 582432 604401
rect 582380 577643 582432 577652
rect 582380 577609 582389 577643
rect 582389 577609 582423 577643
rect 582423 577609 582432 577643
rect 582380 577600 582432 577609
rect 582380 575467 582432 575476
rect 582380 575433 582389 575467
rect 582389 575433 582423 575467
rect 582423 575433 582432 575467
rect 582380 575424 582432 575433
rect 582380 564315 582432 564324
rect 582380 564281 582389 564315
rect 582389 564281 582423 564315
rect 582423 564281 582432 564315
rect 582380 564272 582432 564281
rect 582380 560235 582432 560244
rect 582380 560201 582389 560235
rect 582389 560201 582423 560235
rect 582423 560201 582432 560235
rect 582380 560192 582432 560201
rect 582380 543779 582432 543788
rect 582380 543745 582389 543779
rect 582389 543745 582423 543779
rect 582423 543745 582432 543779
rect 582380 543736 582432 543745
rect 582380 537863 582432 537872
rect 582380 537829 582389 537863
rect 582389 537829 582423 537863
rect 582423 537829 582432 537863
rect 582380 537820 582432 537829
rect 582380 529975 582432 529984
rect 582380 529941 582389 529975
rect 582389 529941 582423 529975
rect 582423 529941 582432 529975
rect 582380 529932 582432 529941
rect 582380 524535 582432 524544
rect 582380 524501 582389 524535
rect 582389 524501 582423 524535
rect 582423 524501 582432 524535
rect 582380 524492 582432 524501
rect 582380 514947 582432 514956
rect 582380 514913 582389 514947
rect 582389 514913 582423 514947
rect 582423 514913 582432 514947
rect 582380 514904 582432 514913
rect 582380 511343 582432 511352
rect 582380 511309 582389 511343
rect 582389 511309 582423 511343
rect 582423 511309 582432 511343
rect 582380 511300 582432 511309
rect 582380 501007 582432 501016
rect 582380 500973 582389 501007
rect 582389 500973 582423 501007
rect 582423 500973 582432 501007
rect 582380 500964 582432 500973
rect 582472 485843 582524 485852
rect 582472 485809 582481 485843
rect 582481 485809 582515 485843
rect 582515 485809 582524 485843
rect 582472 485800 582524 485809
rect 582380 484687 582432 484696
rect 582380 484653 582389 484687
rect 582389 484653 582423 484687
rect 582423 484653 582432 484687
rect 582380 484644 582432 484653
rect 582472 471495 582524 471504
rect 582472 471461 582481 471495
rect 582481 471461 582515 471495
rect 582515 471461 582524 471495
rect 582472 471452 582524 471461
rect 582564 470815 582616 470824
rect 582564 470781 582573 470815
rect 582573 470781 582607 470815
rect 582607 470781 582616 470815
rect 582564 470772 582616 470781
rect 582564 458167 582616 458176
rect 582564 458133 582573 458167
rect 582573 458133 582607 458167
rect 582607 458133 582616 458167
rect 582564 458124 582616 458133
rect 582380 456807 582432 456816
rect 582380 456773 582389 456807
rect 582389 456773 582423 456807
rect 582423 456773 582432 456807
rect 582380 456764 582432 456773
rect 582472 442051 582524 442060
rect 582472 442017 582481 442051
rect 582481 442017 582515 442051
rect 582515 442017 582524 442051
rect 582472 442008 582524 442017
rect 582380 431647 582432 431656
rect 582380 431613 582389 431647
rect 582389 431613 582423 431647
rect 582423 431613 582432 431647
rect 582380 431604 582432 431613
rect 582564 426479 582616 426488
rect 582564 426445 582573 426479
rect 582573 426445 582607 426479
rect 582607 426445 582616 426479
rect 582564 426436 582616 426445
rect 582472 418319 582524 418328
rect 582472 418285 582481 418319
rect 582481 418285 582515 418319
rect 582515 418285 582524 418319
rect 582472 418276 582524 418285
rect 582380 412811 582432 412820
rect 582380 412777 582389 412811
rect 582389 412777 582423 412811
rect 582423 412777 582432 412811
rect 582380 412768 582432 412777
rect 582564 404991 582616 405000
rect 582564 404957 582573 404991
rect 582573 404957 582607 404991
rect 582607 404957 582616 404991
rect 582564 404948 582616 404957
rect 582472 397511 582524 397520
rect 582472 397477 582481 397511
rect 582481 397477 582515 397511
rect 582515 397477 582524 397511
rect 582472 397468 582524 397477
rect 582564 383707 582616 383716
rect 582564 383673 582573 383707
rect 582573 383673 582607 383707
rect 582607 383673 582616 383707
rect 582564 383664 582616 383673
rect 582380 378471 582432 378480
rect 582380 378437 582389 378471
rect 582389 378437 582423 378471
rect 582423 378437 582432 378471
rect 582380 378428 582432 378437
rect 582380 368543 582432 368552
rect 582380 368509 582389 368543
rect 582389 368509 582423 368543
rect 582423 368509 582432 368543
rect 582380 368500 582432 368509
rect 582472 365143 582524 365152
rect 582472 365109 582481 365143
rect 582481 365109 582515 365143
rect 582515 365109 582524 365143
rect 582472 365100 582524 365109
rect 582656 353311 582708 353320
rect 582656 353277 582665 353311
rect 582665 353277 582699 353311
rect 582699 353277 582708 353311
rect 582656 353268 582708 353277
rect 582564 351951 582616 351960
rect 582564 351917 582573 351951
rect 582573 351917 582607 351951
rect 582607 351917 582616 351951
rect 582564 351908 582616 351917
rect 582564 339507 582616 339516
rect 582564 339473 582573 339507
rect 582573 339473 582607 339507
rect 582607 339473 582616 339507
rect 582564 339464 582616 339473
rect 582380 325295 582432 325304
rect 582380 325261 582389 325295
rect 582389 325261 582423 325295
rect 582423 325261 582432 325295
rect 582380 325252 582432 325261
rect 582472 324343 582524 324352
rect 582472 324309 582481 324343
rect 582481 324309 582515 324343
rect 582515 324309 582524 324343
rect 582472 324300 582524 324309
rect 582656 312103 582708 312112
rect 582656 312069 582665 312103
rect 582665 312069 582699 312103
rect 582699 312069 582708 312103
rect 582656 312060 582708 312069
rect 582380 310539 582432 310548
rect 582380 310505 582389 310539
rect 582389 310505 582423 310539
rect 582423 310505 582432 310539
rect 582380 310496 582432 310505
rect 582564 298775 582616 298784
rect 582564 298741 582573 298775
rect 582573 298741 582607 298775
rect 582607 298741 582616 298775
rect 582564 298732 582616 298741
rect 582564 295375 582616 295384
rect 582564 295341 582573 295375
rect 582573 295341 582607 295375
rect 582607 295341 582616 295375
rect 582564 295332 582616 295341
rect 582656 280211 582708 280220
rect 582656 280177 582665 280211
rect 582665 280177 582699 280211
rect 582699 280177 582708 280211
rect 582656 280168 582708 280177
rect 582472 272255 582524 272264
rect 582472 272221 582481 272255
rect 582481 272221 582515 272255
rect 582515 272221 582524 272255
rect 582472 272212 582524 272221
rect 582472 266407 582524 266416
rect 582472 266373 582481 266407
rect 582481 266373 582515 266407
rect 582515 266373 582524 266407
rect 582472 266364 582524 266373
rect 582380 258927 582432 258936
rect 582380 258893 582389 258927
rect 582389 258893 582423 258927
rect 582423 258893 582432 258927
rect 582380 258884 582432 258893
rect 582380 251243 582432 251252
rect 582380 251209 582389 251243
rect 582389 251209 582423 251243
rect 582423 251209 582432 251243
rect 582380 251200 582432 251209
rect 582564 245599 582616 245608
rect 582564 245565 582573 245599
rect 582573 245565 582607 245599
rect 582607 245565 582616 245599
rect 582564 245556 582616 245565
rect 582748 236011 582800 236020
rect 582748 235977 582757 236011
rect 582757 235977 582791 236011
rect 582791 235977 582800 236011
rect 582748 235968 582800 235977
rect 582656 232407 582708 232416
rect 582656 232373 582665 232407
rect 582665 232373 582699 232407
rect 582699 232373 582708 232407
rect 582656 232364 582708 232373
rect 582656 222207 582708 222216
rect 582656 222173 582665 222207
rect 582665 222173 582699 222207
rect 582699 222173 582708 222207
rect 582656 222164 582708 222173
rect 582472 219079 582524 219088
rect 582472 219045 582481 219079
rect 582481 219045 582515 219079
rect 582515 219045 582524 219079
rect 582472 219036 582524 219045
rect 582840 207043 582892 207052
rect 582840 207009 582849 207043
rect 582849 207009 582883 207043
rect 582883 207009 582892 207043
rect 582840 207000 582892 207009
rect 582380 205751 582432 205760
rect 582380 205717 582389 205751
rect 582389 205717 582423 205751
rect 582423 205717 582432 205751
rect 582380 205708 582432 205717
rect 582564 193239 582616 193248
rect 582564 193205 582573 193239
rect 582573 193205 582607 193239
rect 582607 193205 582616 193239
rect 582564 193196 582616 193205
rect 582748 192559 582800 192568
rect 582748 192525 582757 192559
rect 582757 192525 582791 192559
rect 582791 192525 582800 192559
rect 582748 192516 582800 192525
rect 582656 179231 582708 179240
rect 582656 179197 582665 179231
rect 582665 179197 582699 179231
rect 582699 179197 582708 179231
rect 582656 179188 582708 179197
rect 582472 178075 582524 178084
rect 582472 178041 582481 178075
rect 582481 178041 582515 178075
rect 582515 178041 582524 178075
rect 582472 178032 582524 178041
rect 582840 165903 582892 165912
rect 582840 165869 582849 165903
rect 582849 165869 582883 165903
rect 582883 165869 582892 165903
rect 582840 165860 582892 165869
rect 582380 162911 582432 162920
rect 582380 162877 582389 162911
rect 582389 162877 582423 162911
rect 582423 162877 582432 162911
rect 582380 162868 582432 162877
rect 582564 152711 582616 152720
rect 582564 152677 582573 152711
rect 582573 152677 582607 152711
rect 582607 152677 582616 152711
rect 582564 152668 582616 152677
rect 582564 149107 582616 149116
rect 582564 149073 582573 149107
rect 582573 149073 582607 149107
rect 582607 149073 582616 149107
rect 582564 149064 582616 149073
rect 582472 139383 582524 139392
rect 582472 139349 582481 139383
rect 582481 139349 582515 139383
rect 582515 139349 582524 139383
rect 582472 139340 582524 139349
rect 582472 133943 582524 133952
rect 582472 133909 582481 133943
rect 582481 133909 582515 133943
rect 582515 133909 582524 133943
rect 582472 133900 582524 133909
rect 582380 126055 582432 126064
rect 582380 126021 582389 126055
rect 582389 126021 582423 126055
rect 582423 126021 582432 126055
rect 582380 126012 582432 126021
rect 582380 118711 582432 118720
rect 582380 118677 582389 118711
rect 582389 118677 582423 118711
rect 582423 118677 582432 118711
rect 582380 118668 582432 118677
rect 582564 112863 582616 112872
rect 582564 112829 582573 112863
rect 582573 112829 582607 112863
rect 582607 112829 582616 112863
rect 582564 112820 582616 112829
rect 582564 104907 582616 104916
rect 582564 104873 582573 104907
rect 582573 104873 582607 104907
rect 582607 104873 582616 104907
rect 582564 104864 582616 104873
rect 582472 99535 582524 99544
rect 582472 99501 582481 99535
rect 582481 99501 582515 99535
rect 582515 99501 582524 99535
rect 582472 99492 582524 99501
rect 582472 89743 582524 89752
rect 582472 89709 582481 89743
rect 582481 89709 582515 89743
rect 582515 89709 582524 89743
rect 582472 89700 582524 89709
rect 582380 86207 582432 86216
rect 582380 86173 582389 86207
rect 582389 86173 582423 86207
rect 582423 86173 582432 86207
rect 582380 86164 582432 86173
rect 582380 75939 582432 75948
rect 582380 75905 582389 75939
rect 582389 75905 582423 75939
rect 582423 75905 582432 75939
rect 582380 75896 582432 75905
rect 582564 73015 582616 73024
rect 582564 72981 582573 73015
rect 582573 72981 582607 73015
rect 582607 72981 582616 73015
rect 582564 72972 582616 72981
rect 582564 60775 582616 60784
rect 582564 60741 582573 60775
rect 582573 60741 582607 60775
rect 582607 60741 582616 60775
rect 582564 60732 582616 60741
rect 582472 59687 582524 59696
rect 582472 59653 582481 59687
rect 582481 59653 582515 59687
rect 582515 59653 582524 59687
rect 582472 59644 582524 59653
rect 582380 46359 582432 46368
rect 582380 46325 582389 46359
rect 582389 46325 582423 46359
rect 582423 46325 582432 46359
rect 582380 46316 582432 46325
rect 582656 46155 582708 46164
rect 582656 46121 582665 46155
rect 582665 46121 582699 46155
rect 582699 46121 582708 46155
rect 582656 46112 582708 46121
rect 582564 33099 582616 33108
rect 582564 33065 582573 33099
rect 582573 33065 582607 33099
rect 582607 33065 582616 33099
rect 582564 33056 582616 33065
rect 582472 31807 582524 31816
rect 582472 31773 582481 31807
rect 582481 31773 582515 31807
rect 582515 31773 582524 31807
rect 582472 31764 582524 31773
rect 303620 29792 303672 29844
rect 304768 29792 304820 29844
rect 318800 29792 318852 29844
rect 319948 29792 320000 29844
rect 333980 29792 334032 29844
rect 335128 29792 335180 29844
rect 349160 29792 349212 29844
rect 350308 29792 350360 29844
rect 379520 29792 379572 29844
rect 380668 29792 380720 29844
rect 425060 29792 425112 29844
rect 426208 29792 426260 29844
rect 440240 29792 440292 29844
rect 441480 29792 441532 29844
rect 470600 29792 470652 29844
rect 471840 29792 471892 29844
rect 500960 29792 501012 29844
rect 502200 29792 502252 29844
rect 561680 29792 561732 29844
rect 562920 29792 562972 29844
rect 1308 27548 1360 27600
rect 6000 27548 6052 27600
rect 26332 27548 26384 27600
rect 29644 27548 29696 27600
rect 36452 27548 36504 27600
rect 39304 27548 39356 27600
rect 41512 27548 41564 27600
rect 43444 27548 43496 27600
rect 46572 27548 46624 27600
rect 47584 27548 47636 27600
rect 51632 27548 51684 27600
rect 52368 27548 52420 27600
rect 56692 27548 56744 27600
rect 57888 27548 57940 27600
rect 58624 27548 58676 27600
rect 122380 27548 122432 27600
rect 124864 27548 124916 27600
rect 127440 27548 127492 27600
rect 162124 27548 162176 27600
rect 162952 27548 163004 27600
rect 166264 27548 166316 27600
rect 168012 27548 168064 27600
rect 190460 27548 190512 27600
rect 193312 27548 193364 27600
rect 313924 27548 313976 27600
rect 314844 27548 314896 27600
rect 454684 27548 454736 27600
rect 456616 27548 456668 27600
rect 53104 27480 53156 27532
rect 132500 27480 132552 27532
rect 66812 27412 66864 27464
rect 69664 27412 69716 27464
rect 81992 27412 82044 27464
rect 83464 27412 83516 27464
rect 97080 27412 97132 27464
rect 101404 27412 101456 27464
rect 102140 27412 102192 27464
rect 114468 27412 114520 27464
rect 365444 27412 365496 27464
rect 68284 27344 68336 27396
rect 107200 27344 107252 27396
rect 107568 27344 107620 27396
rect 375564 27344 375616 27396
rect 71872 27276 71924 27328
rect 90364 27276 90416 27328
rect 93768 27276 93820 27328
rect 395804 27276 395856 27328
rect 75184 27208 75236 27260
rect 86776 27208 86828 27260
rect 405924 27208 405976 27260
rect 31392 27140 31444 27192
rect 50344 27140 50396 27192
rect 82728 27140 82780 27192
rect 410984 27140 411036 27192
rect 486424 27140 486476 27192
rect 33784 27072 33836 27124
rect 486976 27072 487028 27124
rect 527456 27072 527508 27124
rect 5448 27004 5500 27056
rect 11060 27004 11112 27056
rect 32404 27004 32456 27056
rect 497096 27004 497148 27056
rect 497464 27004 497516 27056
rect 517336 27004 517388 27056
rect 518164 27004 518216 27056
rect 532516 27004 532568 27056
rect 4068 26936 4120 26988
rect 16120 26936 16172 26988
rect 36544 26936 36596 26988
rect 567936 26936 567988 26988
rect 6828 26868 6880 26920
rect 21180 26868 21232 26920
rect 35164 26868 35216 26920
rect 578148 26868 578200 26920
rect 65524 26800 65576 26852
rect 117320 26800 117372 26852
rect 79324 26732 79376 26784
rect 92020 26732 92072 26784
rect 40684 25712 40736 25764
rect 157340 25712 157392 25764
rect 18604 25644 18656 25696
rect 182180 25644 182232 25696
rect 54484 25576 54536 25628
rect 451280 25576 451332 25628
rect 7564 25508 7616 25560
rect 552020 25508 552072 25560
rect 11704 24080 11756 24132
rect 506480 24080 506532 24132
rect 119988 22720 120040 22772
rect 190460 22720 190512 22772
rect 29644 21360 29696 21412
rect 122840 21360 122892 21412
rect 25504 19932 25556 19984
rect 172520 19932 172572 19984
rect 582656 19839 582708 19848
rect 582656 19805 582665 19839
rect 582665 19805 582699 19839
rect 582699 19805 582708 19839
rect 582656 19796 582708 19805
rect 62028 18572 62080 18624
rect 98000 18572 98052 18624
rect 52368 17212 52420 17264
rect 104900 17212 104952 17264
rect 69664 15920 69716 15972
rect 94688 15920 94740 15972
rect 51724 15852 51776 15904
rect 142160 15852 142212 15904
rect 144736 15852 144788 15904
rect 536840 15852 536892 15904
rect 41328 14424 41380 14476
rect 303620 14424 303672 14476
rect 22744 13064 22796 13116
rect 178040 13064 178092 13116
rect 70308 11772 70360 11824
rect 101404 11772 101456 11824
rect 39304 11704 39356 11756
rect 116400 11704 116452 11756
rect 125876 11704 125928 11756
rect 486424 11704 486476 11756
rect 39304 10344 39356 10396
rect 151820 10344 151872 10396
rect 14464 10276 14516 10328
rect 557540 10276 557592 10328
rect 27712 9120 27764 9172
rect 162124 9120 162176 9172
rect 44272 9052 44324 9104
rect 299480 9052 299532 9104
rect 49884 8984 49936 9036
rect 136640 8984 136692 9036
rect 141240 8984 141292 9036
rect 542360 8984 542412 9036
rect 50160 8916 50212 8968
rect 454684 8916 454736 8968
rect 122288 7964 122340 8016
rect 187700 7964 187752 8016
rect 23020 7896 23072 7948
rect 166264 7896 166316 7948
rect 37188 7828 37240 7880
rect 309140 7828 309192 7880
rect 33600 7760 33652 7812
rect 313924 7760 313976 7812
rect 50344 7692 50396 7744
rect 119896 7692 119948 7744
rect 132960 7692 133012 7744
rect 497464 7692 497516 7744
rect 43168 7624 43220 7676
rect 147680 7624 147732 7676
rect 148324 7624 148376 7676
rect 518164 7624 518216 7676
rect 43444 7556 43496 7608
rect 112812 7556 112864 7608
rect 129372 7556 129424 7608
rect 521660 7556 521712 7608
rect 80888 6808 80940 6860
rect 86960 6808 87012 6860
rect 77208 6672 77260 6724
rect 87972 6672 88024 6724
rect 63224 6604 63276 6656
rect 111800 6604 111852 6656
rect 115204 6604 115256 6656
rect 197360 6604 197412 6656
rect 582472 6647 582524 6656
rect 582472 6613 582481 6647
rect 582481 6613 582515 6647
rect 582515 6613 582524 6647
rect 582472 6604 582524 6613
rect 47584 6536 47636 6588
rect 109316 6536 109368 6588
rect 111616 6536 111668 6588
rect 202880 6536 202932 6588
rect 57888 6468 57940 6520
rect 102232 6468 102284 6520
rect 108120 6468 108172 6520
rect 208400 6468 208452 6520
rect 30104 6400 30156 6452
rect 318800 6400 318852 6452
rect 26516 6332 26568 6384
rect 324320 6332 324372 6384
rect 21824 6264 21876 6316
rect 329840 6264 329892 6316
rect 17040 6196 17092 6248
rect 333980 6196 334032 6248
rect 52552 6128 52604 6180
rect 124864 6128 124916 6180
rect 136456 6128 136508 6180
rect 512000 6128 512052 6180
rect 76196 5448 76248 5500
rect 253940 5448 253992 5500
rect 72608 5380 72660 5432
rect 258080 5380 258132 5432
rect 69112 5312 69164 5364
rect 263600 5312 263652 5364
rect 65616 5244 65668 5296
rect 269120 5244 269172 5296
rect 62028 5176 62080 5228
rect 273260 5176 273312 5228
rect 58440 5108 58492 5160
rect 278780 5108 278832 5160
rect 54944 5040 54996 5092
rect 284300 5040 284352 5092
rect 51356 4972 51408 5024
rect 288440 4972 288492 5024
rect 47860 4904 47912 4956
rect 293960 4904 294012 4956
rect 12348 4836 12400 4888
rect 339500 4836 339552 4888
rect 7656 4768 7708 4820
rect 345020 4768 345072 4820
rect 73804 4700 73856 4752
rect 75184 4700 75236 4752
rect 83464 4700 83516 4752
rect 84476 4700 84528 4752
rect 79692 4564 79744 4616
rect 248420 4700 248472 4752
rect 83280 4496 83332 4548
rect 242900 4632 242952 4684
rect 86868 4428 86920 4480
rect 238760 4564 238812 4616
rect 90456 4496 90508 4548
rect 233240 4496 233292 4548
rect 93952 4428 94004 4480
rect 227720 4428 227772 4480
rect 59636 4360 59688 4412
rect 65524 4360 65576 4412
rect 97448 4360 97500 4412
rect 223580 4360 223632 4412
rect 101036 4292 101088 4344
rect 218060 4292 218112 4344
rect 104532 4224 104584 4276
rect 212540 4224 212592 4276
rect 48964 4156 49016 4208
rect 53104 4156 53156 4208
rect 56048 4156 56100 4208
rect 58624 4156 58676 4208
rect 66720 4156 66772 4208
rect 68284 4156 68336 4208
rect 77392 4156 77444 4208
rect 79324 4156 79376 4208
rect 90364 4156 90416 4208
rect 91560 4156 91612 4208
rect 1676 4088 1728 4140
rect 7564 4088 7616 4140
rect 75000 4088 75052 4140
rect 420920 4088 420972 4140
rect 71504 4020 71556 4072
rect 425060 4020 425112 4072
rect 67916 3952 67968 4004
rect 430580 3952 430632 4004
rect 64328 3884 64380 3936
rect 436100 3884 436152 3936
rect 45468 3816 45520 3868
rect 49884 3816 49936 3868
rect 60832 3816 60884 3868
rect 440240 3816 440292 3868
rect 41880 3748 41932 3800
rect 51724 3748 51776 3800
rect 57244 3748 57296 3800
rect 445760 3748 445812 3800
rect 13544 3680 13596 3732
rect 22744 3680 22796 3732
rect 31300 3680 31352 3732
rect 40684 3680 40736 3732
rect 46664 3680 46716 3732
rect 460940 3680 460992 3732
rect 19432 3612 19484 3664
rect 32404 3612 32456 3664
rect 34796 3612 34848 3664
rect 39304 3612 39356 3664
rect 43076 3612 43128 3664
rect 466460 3612 466512 3664
rect 8760 3544 8812 3596
rect 18604 3544 18656 3596
rect 20628 3544 20680 3596
rect 36544 3544 36596 3596
rect 39580 3544 39632 3596
rect 470600 3544 470652 3596
rect 572 3476 624 3528
rect 1308 3476 1360 3528
rect 11152 3476 11204 3528
rect 2872 3408 2924 3460
rect 14464 3408 14516 3460
rect 28908 3476 28960 3528
rect 33784 3476 33836 3528
rect 40684 3476 40736 3528
rect 41328 3476 41380 3528
rect 35164 3408 35216 3460
rect 35992 3340 36044 3392
rect 476120 3476 476172 3528
rect 53748 3408 53800 3460
rect 54484 3408 54536 3460
rect 38384 3272 38436 3324
rect 43168 3272 43220 3324
rect 32404 3204 32456 3256
rect 481640 3408 481692 3460
rect 547788 3408 547840 3460
rect 579804 3408 579856 3460
rect 82084 3340 82136 3392
rect 82728 3340 82780 3392
rect 85672 3340 85724 3392
rect 86776 3340 86828 3392
rect 78588 3272 78640 3324
rect 415400 3340 415452 3392
rect 92756 3272 92808 3324
rect 93768 3272 93820 3324
rect 89168 3204 89220 3256
rect 400220 3272 400272 3324
rect 96252 3136 96304 3188
rect 390560 3204 390612 3256
rect 99840 3136 99892 3188
rect 385040 3136 385092 3188
rect 18236 3068 18288 3120
rect 25504 3068 25556 3120
rect 103336 3068 103388 3120
rect 379520 3068 379572 3120
rect 106924 3000 106976 3052
rect 107568 3000 107620 3052
rect 110512 3000 110564 3052
rect 369860 3000 369912 3052
rect 9956 2932 10008 2984
rect 11704 2932 11756 2984
rect 114008 2932 114060 2984
rect 114468 2932 114520 2984
rect 118792 2932 118844 2984
rect 119988 2932 120040 2984
rect 117596 2864 117648 2916
rect 360200 2932 360252 2984
rect 121092 2864 121144 2916
rect 354680 2864 354732 2916
rect 124680 2796 124732 2848
rect 349160 2796 349212 2848
<< metal2 >>
rect 6932 703582 7972 703610
rect 18 683768 74 683777
rect 18 683703 74 683712
rect 32 645425 60 683703
rect 6932 681698 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 89364 703582 89668 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 24320 699718 24348 703520
rect 40512 700398 40540 703520
rect 72988 703050 73016 703520
rect 89180 703474 89208 703520
rect 89364 703474 89392 703582
rect 89180 703446 89392 703474
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 41328 700334 41380 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 24780 681698 24808 699654
rect 6092 681692 6144 681698
rect 6092 681634 6144 681640
rect 6920 681692 6972 681698
rect 6920 681634 6972 681640
rect 24768 681692 24820 681698
rect 24768 681634 24820 681640
rect 27988 681692 28040 681698
rect 27988 681634 28040 681640
rect 6104 678858 6132 681634
rect 6056 678830 6132 678858
rect 28000 678858 28028 681634
rect 41340 681018 41368 700334
rect 41328 681012 41380 681018
rect 41328 680954 41380 680960
rect 49976 681012 50028 681018
rect 49976 680954 50028 680960
rect 49988 678858 50016 680954
rect 71792 678858 71820 702986
rect 89640 681698 89668 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 154316 703582 154528 703610
rect 105464 700398 105492 703520
rect 137848 702434 137876 703520
rect 154132 703474 154160 703520
rect 154316 703474 154344 703582
rect 154132 703446 154344 703474
rect 137848 702406 137968 702434
rect 105452 700392 105504 700398
rect 105452 700334 105504 700340
rect 106188 700392 106240 700398
rect 106188 700334 106240 700340
rect 89628 681692 89680 681698
rect 89628 681634 89680 681640
rect 93952 681692 94004 681698
rect 93952 681634 94004 681640
rect 93964 678858 93992 681634
rect 106200 681018 106228 700334
rect 106188 681012 106240 681018
rect 106188 680954 106240 680960
rect 115940 681012 115992 681018
rect 115940 680954 115992 680960
rect 115952 678858 115980 680954
rect 137940 680354 137968 702406
rect 154500 680678 154528 703582
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 284036 703582 284248 703610
rect 170324 700262 170352 703520
rect 170312 700256 170364 700262
rect 170312 700198 170364 700204
rect 171048 700256 171100 700262
rect 171048 700198 171100 700204
rect 171060 681018 171088 700198
rect 171048 681012 171100 681018
rect 171048 680954 171100 680960
rect 181996 681012 182048 681018
rect 181996 680954 182048 680960
rect 154488 680672 154540 680678
rect 154488 680614 154540 680620
rect 160008 680672 160060 680678
rect 160008 680614 160060 680620
rect 137940 680326 138060 680354
rect 138032 678994 138060 680326
rect 138032 678966 138104 678994
rect 28000 678830 28072 678858
rect 49988 678830 50060 678858
rect 71792 678830 72048 678858
rect 93964 678830 94036 678858
rect 115952 678830 116024 678858
rect 6056 678776 6084 678830
rect 28044 678776 28072 678830
rect 50032 678776 50060 678830
rect 72020 678776 72048 678830
rect 94008 678776 94036 678830
rect 115996 678776 116024 678830
rect 138076 678776 138104 678966
rect 160020 678858 160048 680614
rect 182008 678858 182036 680954
rect 202800 680950 202828 703520
rect 218992 702434 219020 703520
rect 218992 702406 219388 702434
rect 219360 681018 219388 702406
rect 235184 700398 235212 703520
rect 235172 700392 235224 700398
rect 235172 700334 235224 700340
rect 235908 700392 235960 700398
rect 235908 700334 235960 700340
rect 235920 681018 235948 700334
rect 267660 681290 267688 703520
rect 283852 703474 283880 703520
rect 284036 703474 284064 703582
rect 283852 703446 284064 703474
rect 267648 681284 267700 681290
rect 267648 681226 267700 681232
rect 270040 681284 270092 681290
rect 270040 681226 270092 681232
rect 219348 681012 219400 681018
rect 219348 680954 219400 680960
rect 225972 681012 226024 681018
rect 225972 680954 226024 680960
rect 235908 681012 235960 681018
rect 235908 680954 235960 680960
rect 248052 681012 248104 681018
rect 248052 680954 248104 680960
rect 202788 680944 202840 680950
rect 202788 680886 202840 680892
rect 203984 680944 204036 680950
rect 203984 680886 204036 680892
rect 203996 678858 204024 680886
rect 225984 678858 226012 680954
rect 248064 678858 248092 680954
rect 270052 678858 270080 681226
rect 284220 681018 284248 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 300136 699718 300164 703520
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 300768 699712 300820 699718
rect 300768 699654 300820 699660
rect 300780 681018 300808 699654
rect 332520 681154 332548 703520
rect 348804 702434 348832 703520
rect 348804 702406 349108 702434
rect 332508 681148 332560 681154
rect 332508 681090 332560 681096
rect 336004 681148 336056 681154
rect 336004 681090 336056 681096
rect 284208 681012 284260 681018
rect 284208 680954 284260 680960
rect 292028 681012 292080 681018
rect 292028 680954 292080 680960
rect 300768 681012 300820 681018
rect 300768 680954 300820 680960
rect 314016 681012 314068 681018
rect 314016 680954 314068 680960
rect 292040 678858 292068 680954
rect 314028 678858 314056 680954
rect 336016 678858 336044 681090
rect 349080 681018 349108 702406
rect 364996 700534 365024 703520
rect 364984 700528 365036 700534
rect 364984 700470 365036 700476
rect 365628 700528 365680 700534
rect 365628 700470 365680 700476
rect 365640 681018 365668 700470
rect 397472 699990 397500 703520
rect 413664 702434 413692 703520
rect 413664 702406 413968 702434
rect 397460 699984 397512 699990
rect 397460 699926 397512 699932
rect 398748 699984 398800 699990
rect 398748 699926 398800 699932
rect 349068 681012 349120 681018
rect 349068 680954 349120 680960
rect 358084 681012 358136 681018
rect 358084 680954 358136 680960
rect 365628 681012 365680 681018
rect 365628 680954 365680 680960
rect 380072 681012 380124 681018
rect 380072 680954 380124 680960
rect 358096 678858 358124 680954
rect 380084 678858 380112 680954
rect 398760 680746 398788 699926
rect 413940 681018 413968 702406
rect 429856 699718 429884 703520
rect 462332 699718 462360 703520
rect 478524 702434 478552 703520
rect 478524 702406 478828 702434
rect 429844 699712 429896 699718
rect 429844 699654 429896 699660
rect 430488 699712 430540 699718
rect 430488 699654 430540 699660
rect 462320 699712 462372 699718
rect 462320 699654 462372 699660
rect 463608 699712 463660 699718
rect 463608 699654 463660 699660
rect 430500 681018 430528 699654
rect 413928 681012 413980 681018
rect 413928 680954 413980 680960
rect 424048 681012 424100 681018
rect 424048 680954 424100 680960
rect 430488 681012 430540 681018
rect 430488 680954 430540 680960
rect 446036 681012 446088 681018
rect 446036 680954 446088 680960
rect 398748 680740 398800 680746
rect 398748 680682 398800 680688
rect 402060 680740 402112 680746
rect 402060 680682 402112 680688
rect 402072 678858 402100 680682
rect 424060 678858 424088 680954
rect 446048 678858 446076 680954
rect 463620 680950 463648 699654
rect 478800 681018 478828 702406
rect 494808 699718 494836 703520
rect 527192 700534 527220 703520
rect 543476 702434 543504 703520
rect 543476 702406 543688 702434
rect 527180 700528 527232 700534
rect 527180 700470 527232 700476
rect 528468 700528 528520 700534
rect 528468 700470 528520 700476
rect 494796 699712 494848 699718
rect 494796 699654 494848 699660
rect 495348 699712 495400 699718
rect 495348 699654 495400 699660
rect 495360 681018 495388 699654
rect 528480 681018 528508 700470
rect 543660 681018 543688 702406
rect 559668 699718 559696 703520
rect 559656 699712 559708 699718
rect 559656 699654 559708 699660
rect 560208 699712 560260 699718
rect 560208 699654 560260 699660
rect 560220 681018 560248 699654
rect 582378 697232 582434 697241
rect 582378 697167 582380 697176
rect 582432 697167 582434 697176
rect 582380 697138 582432 697144
rect 582470 683904 582526 683913
rect 582470 683839 582472 683848
rect 582524 683839 582526 683848
rect 582472 683810 582524 683816
rect 478788 681012 478840 681018
rect 478788 680954 478840 680960
rect 490104 681012 490156 681018
rect 490104 680954 490156 680960
rect 495348 681012 495400 681018
rect 495348 680954 495400 680960
rect 512092 681012 512144 681018
rect 512092 680954 512144 680960
rect 528468 681012 528520 681018
rect 528468 680954 528520 680960
rect 534080 681012 534132 681018
rect 534080 680954 534132 680960
rect 543648 681012 543700 681018
rect 543648 680954 543700 680960
rect 556068 681012 556120 681018
rect 556068 680954 556120 680960
rect 560208 681012 560260 681018
rect 560208 680954 560260 680960
rect 578056 681012 578108 681018
rect 578056 680954 578108 680960
rect 463608 680944 463660 680950
rect 463608 680886 463660 680892
rect 468116 680944 468168 680950
rect 468116 680886 468168 680892
rect 468128 678858 468156 680886
rect 490116 678858 490144 680954
rect 512104 678858 512132 680954
rect 534092 678858 534120 680954
rect 556080 678858 556108 680954
rect 578068 678858 578096 680954
rect 160020 678830 160092 678858
rect 182008 678830 182080 678858
rect 203996 678830 204068 678858
rect 225984 678830 226056 678858
rect 248064 678830 248136 678858
rect 270052 678830 270124 678858
rect 292040 678830 292112 678858
rect 314028 678830 314100 678858
rect 336016 678830 336088 678858
rect 358096 678830 358168 678858
rect 380084 678830 380156 678858
rect 402072 678830 402144 678858
rect 424060 678830 424132 678858
rect 446048 678830 446120 678858
rect 468128 678830 468200 678858
rect 490116 678830 490188 678858
rect 512104 678830 512176 678858
rect 534092 678830 534164 678858
rect 556080 678830 556152 678858
rect 578068 678830 578140 678858
rect 160064 678776 160092 678830
rect 182052 678776 182080 678830
rect 204040 678776 204068 678830
rect 226028 678776 226056 678830
rect 248108 678776 248136 678830
rect 270096 678776 270124 678830
rect 292084 678776 292112 678830
rect 314072 678776 314100 678830
rect 336060 678776 336088 678830
rect 358140 678776 358168 678830
rect 380128 678776 380156 678830
rect 402116 678776 402144 678830
rect 424104 678776 424132 678830
rect 446092 678776 446120 678830
rect 468172 678776 468200 678830
rect 490160 678776 490188 678830
rect 512148 678776 512176 678830
rect 534136 678776 534164 678830
rect 556124 678776 556152 678830
rect 578112 678776 578140 678830
rect 582380 677544 582432 677550
rect 582380 677486 582432 677492
rect 582392 676841 582420 677486
rect 110 676832 166 676841
rect 110 676767 166 676776
rect 582378 676832 582434 676841
rect 582378 676767 582434 676776
rect 124 658238 152 676767
rect 2778 671256 2834 671265
rect 2778 671191 2834 671200
rect 2792 661201 2820 671191
rect 582380 670744 582432 670750
rect 582378 670712 582380 670721
rect 582432 670712 582434 670721
rect 582378 670647 582434 670656
rect 582472 662380 582524 662386
rect 582472 662322 582524 662328
rect 582484 662153 582512 662322
rect 582470 662144 582526 662153
rect 582470 662079 582526 662088
rect 2778 661192 2834 661201
rect 2778 661127 2834 661136
rect 112 658232 164 658238
rect 572 658232 624 658238
rect 112 658174 164 658180
rect 570 658200 572 658209
rect 624 658200 626 658209
rect 570 658135 626 658144
rect 582380 648576 582432 648582
rect 582380 648518 582432 648524
rect 582392 647601 582420 648518
rect 582378 647592 582434 647601
rect 582378 647527 582434 647536
rect 18 645416 74 645425
rect 18 645351 74 645360
rect 582378 644056 582434 644065
rect 582378 643991 582380 644000
rect 582432 643991 582434 644000
rect 582380 643962 582432 643968
rect 582380 633412 582432 633418
rect 582380 633354 582432 633360
rect 582392 632913 582420 633354
rect 582378 632904 582434 632913
rect 582378 632839 582434 632848
rect 20 632120 72 632126
rect 572 632120 624 632126
rect 20 632062 72 632068
rect 570 632088 572 632097
rect 624 632088 626 632097
rect 32 598233 60 632062
rect 570 632023 626 632032
rect 582378 630864 582434 630873
rect 582378 630799 582380 630808
rect 582432 630799 582434 630808
rect 582380 630770 582432 630776
rect 110 629640 166 629649
rect 110 629575 166 629584
rect 124 606665 152 629575
rect 202 618624 258 618633
rect 202 618559 258 618568
rect 216 614009 244 618559
rect 582380 618248 582432 618254
rect 582378 618216 582380 618225
rect 582432 618216 582434 618225
rect 582378 618151 582434 618160
rect 582378 617536 582434 617545
rect 582378 617471 582380 617480
rect 582432 617471 582434 617480
rect 582380 617442 582432 617448
rect 202 614000 258 614009
rect 202 613935 258 613944
rect 110 606656 166 606665
rect 110 606591 166 606600
rect 582380 604444 582432 604450
rect 582380 604386 582432 604392
rect 582392 603673 582420 604386
rect 582378 603664 582434 603673
rect 582378 603599 582434 603608
rect 18 598224 74 598233
rect 18 598159 74 598168
rect 580722 591016 580778 591025
rect 580722 590951 580778 590960
rect 580736 588973 580764 590951
rect 580722 588964 580778 588973
rect 580722 588899 580778 588908
rect 110 582448 166 582457
rect 110 582383 166 582392
rect 18 579728 74 579737
rect 18 579663 74 579672
rect 32 551041 60 579663
rect 124 554441 152 582383
rect 582378 577688 582434 577697
rect 582378 577623 582380 577632
rect 582432 577623 582434 577632
rect 582380 577594 582432 577600
rect 582380 575476 582432 575482
rect 582380 575418 582432 575424
rect 582392 574297 582420 575418
rect 582378 574288 582434 574297
rect 582378 574223 582434 574232
rect 582378 564360 582434 564369
rect 582378 564295 582380 564304
rect 582432 564295 582434 564304
rect 582380 564266 582432 564272
rect 582380 560244 582432 560250
rect 582380 560186 582432 560192
rect 582392 559745 582420 560186
rect 582378 559736 582434 559745
rect 582378 559671 582434 559680
rect 110 554432 166 554441
rect 110 554367 166 554376
rect 18 551032 74 551041
rect 18 550967 74 550976
rect 582378 544912 582434 544921
rect 582378 544847 582434 544856
rect 582392 543794 582420 544847
rect 582380 543788 582432 543794
rect 582380 543730 582432 543736
rect 582380 537872 582432 537878
rect 582378 537840 582380 537849
rect 582432 537840 582434 537849
rect 582378 537775 582434 537784
rect 18 535256 74 535265
rect 18 535191 74 535200
rect 32 502353 60 535191
rect 582378 530224 582434 530233
rect 582378 530159 582434 530168
rect 582392 529990 582420 530159
rect 582380 529984 582432 529990
rect 582380 529926 582432 529932
rect 110 527368 166 527377
rect 110 527303 166 527312
rect 124 503985 152 527303
rect 582380 524544 582432 524550
rect 582378 524512 582380 524521
rect 582432 524512 582434 524521
rect 582378 524447 582434 524456
rect 2686 519480 2742 519489
rect 2686 519415 2742 519424
rect 2700 514865 2728 519415
rect 582378 515672 582434 515681
rect 582378 515607 582434 515616
rect 582392 514962 582420 515607
rect 582380 514956 582432 514962
rect 582380 514898 582432 514904
rect 2686 514856 2742 514865
rect 2686 514791 2742 514800
rect 582380 511352 582432 511358
rect 582378 511320 582380 511329
rect 582432 511320 582434 511329
rect 582378 511255 582434 511264
rect 110 503976 166 503985
rect 110 503911 166 503920
rect 18 502344 74 502353
rect 18 502279 74 502288
rect 582380 501016 582432 501022
rect 582378 500984 582380 500993
rect 582432 500984 582434 500993
rect 582378 500919 582434 500928
rect 18 488200 74 488209
rect 18 488135 74 488144
rect 32 449857 60 488135
rect 582470 486296 582526 486305
rect 582470 486231 582526 486240
rect 582484 485858 582512 486231
rect 582472 485852 582524 485858
rect 582472 485794 582524 485800
rect 582380 484696 582432 484702
rect 582378 484664 582380 484673
rect 582432 484664 582434 484673
rect 582378 484599 582434 484608
rect 110 475144 166 475153
rect 110 475079 166 475088
rect 124 456793 152 475079
rect 2778 472424 2834 472433
rect 2778 472359 2834 472368
rect 2792 462641 2820 472359
rect 582562 471744 582618 471753
rect 582562 471679 582618 471688
rect 582472 471504 582524 471510
rect 582470 471472 582472 471481
rect 582524 471472 582526 471481
rect 582470 471407 582526 471416
rect 582576 470830 582604 471679
rect 582564 470824 582616 470830
rect 582564 470766 582616 470772
rect 2778 462632 2834 462641
rect 2778 462567 2834 462576
rect 582564 458176 582616 458182
rect 582562 458144 582564 458153
rect 582616 458144 582618 458153
rect 582562 458079 582618 458088
rect 582378 457056 582434 457065
rect 582378 456991 582434 457000
rect 582392 456822 582420 456991
rect 582380 456816 582432 456822
rect 110 456784 166 456793
rect 582380 456758 582432 456764
rect 110 456719 166 456728
rect 18 449848 74 449857
rect 18 449783 74 449792
rect 582470 442368 582526 442377
rect 582470 442303 582526 442312
rect 582484 442066 582512 442303
rect 582472 442060 582524 442066
rect 582472 442002 582524 442008
rect 18 441008 74 441017
rect 18 440943 74 440952
rect 32 398041 60 440943
rect 582380 431656 582432 431662
rect 582378 431624 582380 431633
rect 582432 431624 582434 431633
rect 582378 431559 582434 431568
rect 582562 427816 582618 427825
rect 582562 427751 582618 427760
rect 582576 426494 582604 427751
rect 582564 426488 582616 426494
rect 582564 426430 582616 426436
rect 110 425232 166 425241
rect 110 425167 166 425176
rect 124 411097 152 425167
rect 2778 423600 2834 423609
rect 2778 423535 2834 423544
rect 110 411088 166 411097
rect 110 411023 166 411032
rect 2792 409465 2820 423535
rect 582472 418328 582524 418334
rect 582470 418296 582472 418305
rect 582524 418296 582526 418305
rect 582470 418231 582526 418240
rect 582378 412992 582434 413001
rect 582378 412927 582434 412936
rect 582392 412826 582420 412927
rect 582380 412820 582432 412826
rect 582380 412762 582432 412768
rect 2778 409456 2834 409465
rect 2778 409391 2834 409400
rect 582564 405000 582616 405006
rect 582562 404968 582564 404977
rect 582616 404968 582618 404977
rect 582562 404903 582618 404912
rect 582470 398440 582526 398449
rect 582470 398375 582526 398384
rect 18 398032 74 398041
rect 18 397967 74 397976
rect 582484 397526 582512 398375
rect 582472 397520 582524 397526
rect 582472 397462 582524 397468
rect 110 393816 166 393825
rect 110 393751 166 393760
rect 18 378040 74 378049
rect 18 377975 74 377984
rect 32 358737 60 377975
rect 18 358728 74 358737
rect 18 358663 74 358672
rect 18 346624 74 346633
rect 18 346559 74 346568
rect 32 293729 60 346559
rect 124 345953 152 393751
rect 582562 383752 582618 383761
rect 582562 383687 582564 383696
rect 582616 383687 582618 383696
rect 582564 383658 582616 383664
rect 582380 378480 582432 378486
rect 582378 378448 582380 378457
rect 582432 378448 582434 378457
rect 582378 378383 582434 378392
rect 2778 371376 2834 371385
rect 2778 371311 2834 371320
rect 2792 362273 2820 371311
rect 582378 369064 582434 369073
rect 582378 368999 582434 369008
rect 582392 368558 582420 368999
rect 582380 368552 582432 368558
rect 582380 368494 582432 368500
rect 582472 365152 582524 365158
rect 582470 365120 582472 365129
rect 582524 365120 582526 365129
rect 582470 365055 582526 365064
rect 2778 362264 2834 362273
rect 2778 362199 2834 362208
rect 582654 354512 582710 354521
rect 582654 354447 582710 354456
rect 582668 353326 582696 354447
rect 582656 353320 582708 353326
rect 582656 353262 582708 353268
rect 582564 351960 582616 351966
rect 582562 351928 582564 351937
rect 582616 351928 582618 351937
rect 582562 351863 582618 351872
rect 110 345944 166 345953
rect 110 345879 166 345888
rect 582562 339824 582618 339833
rect 582562 339759 582618 339768
rect 582576 339522 582604 339759
rect 582564 339516 582616 339522
rect 582564 339458 582616 339464
rect 110 330984 166 330993
rect 110 330919 166 330928
rect 124 306513 152 330919
rect 582380 325304 582432 325310
rect 582378 325272 582380 325281
rect 582432 325272 582434 325281
rect 582378 325207 582434 325216
rect 582470 325136 582526 325145
rect 582470 325071 582526 325080
rect 582484 324358 582512 325071
rect 582472 324352 582524 324358
rect 582472 324294 582524 324300
rect 2778 319288 2834 319297
rect 2778 319223 2834 319232
rect 2792 315217 2820 319223
rect 2778 315208 2834 315217
rect 2778 315143 2834 315152
rect 582656 312112 582708 312118
rect 582654 312080 582656 312089
rect 582708 312080 582710 312089
rect 582654 312015 582710 312024
rect 582378 310584 582434 310593
rect 582378 310519 582380 310528
rect 582432 310519 582434 310528
rect 582380 310490 582432 310496
rect 110 306504 166 306513
rect 110 306439 166 306448
rect 110 299432 166 299441
rect 110 299367 166 299376
rect 18 293720 74 293729
rect 18 293655 74 293664
rect 18 283656 74 283665
rect 18 283591 74 283600
rect 32 254697 60 283591
rect 18 254688 74 254697
rect 18 254623 74 254632
rect 18 252240 74 252249
rect 18 252175 74 252184
rect 32 189145 60 252175
rect 124 241505 152 299367
rect 582564 298784 582616 298790
rect 582562 298752 582564 298761
rect 582616 298752 582618 298761
rect 582562 298687 582618 298696
rect 582562 295896 582618 295905
rect 582562 295831 582618 295840
rect 582576 295390 582604 295831
rect 582564 295384 582616 295390
rect 582564 295326 582616 295332
rect 582654 281072 582710 281081
rect 582654 281007 582710 281016
rect 582668 280226 582696 281007
rect 582656 280220 582708 280226
rect 582656 280162 582708 280168
rect 582472 272264 582524 272270
rect 582470 272232 582472 272241
rect 582524 272232 582526 272241
rect 582470 272167 582526 272176
rect 582470 266520 582526 266529
rect 582470 266455 582526 266464
rect 582484 266422 582512 266455
rect 582472 266416 582524 266422
rect 582472 266358 582524 266364
rect 582380 258936 582432 258942
rect 582378 258904 582380 258913
rect 582432 258904 582434 258913
rect 582378 258839 582434 258848
rect 582378 251832 582434 251841
rect 582378 251767 582434 251776
rect 582392 251258 582420 251767
rect 582380 251252 582432 251258
rect 582380 251194 582432 251200
rect 582564 245608 582616 245614
rect 582562 245576 582564 245585
rect 582616 245576 582618 245585
rect 582562 245511 582618 245520
rect 110 241496 166 241505
rect 110 241431 166 241440
rect 582746 237280 582802 237289
rect 582746 237215 582802 237224
rect 110 236464 166 236473
rect 110 236399 166 236408
rect 124 202473 152 236399
rect 582760 236026 582788 237215
rect 582748 236020 582800 236026
rect 582748 235962 582800 235968
rect 582656 232416 582708 232422
rect 582654 232384 582656 232393
rect 582708 232384 582710 232393
rect 582654 232319 582710 232328
rect 582654 222592 582710 222601
rect 582654 222527 582710 222536
rect 582668 222222 582696 222527
rect 582656 222216 582708 222222
rect 582656 222158 582708 222164
rect 2042 220824 2098 220833
rect 2042 220759 2098 220768
rect 2056 214985 2084 220759
rect 582472 219088 582524 219094
rect 582470 219056 582472 219065
rect 582524 219056 582526 219065
rect 582470 218991 582526 219000
rect 2042 214976 2098 214985
rect 2042 214911 2098 214920
rect 582838 207904 582894 207913
rect 582838 207839 582894 207848
rect 582852 207058 582880 207839
rect 582840 207052 582892 207058
rect 582840 206994 582892 207000
rect 582380 205760 582432 205766
rect 582378 205728 582380 205737
rect 582432 205728 582434 205737
rect 582378 205663 582434 205672
rect 2042 205048 2098 205057
rect 2042 204983 2098 204992
rect 110 202464 166 202473
rect 110 202399 166 202408
rect 110 189408 166 189417
rect 110 189343 166 189352
rect 18 189136 74 189145
rect 18 189071 74 189080
rect 18 157992 74 158001
rect 18 157927 74 157936
rect 32 85241 60 157927
rect 124 150385 152 189343
rect 110 150376 166 150385
rect 110 150311 166 150320
rect 2056 136785 2084 204983
rect 582562 193352 582618 193361
rect 582562 193287 582618 193296
rect 582576 193254 582604 193287
rect 582564 193248 582616 193254
rect 582564 193190 582616 193196
rect 582748 192568 582800 192574
rect 582746 192536 582748 192545
rect 582800 192536 582802 192545
rect 582746 192471 582802 192480
rect 582656 179240 582708 179246
rect 582654 179208 582656 179217
rect 582708 179208 582710 179217
rect 582654 179143 582710 179152
rect 582470 178664 582526 178673
rect 582470 178599 582526 178608
rect 582484 178090 582512 178599
rect 582472 178084 582524 178090
rect 582472 178026 582524 178032
rect 2778 173632 2834 173641
rect 2778 173567 2834 173576
rect 2792 162897 2820 173567
rect 582840 165912 582892 165918
rect 582838 165880 582840 165889
rect 582892 165880 582894 165889
rect 582838 165815 582894 165824
rect 582378 163976 582434 163985
rect 582378 163911 582434 163920
rect 582392 162926 582420 163911
rect 582380 162920 582432 162926
rect 2778 162888 2834 162897
rect 582380 162862 582432 162868
rect 2778 162823 2834 162832
rect 582564 152720 582616 152726
rect 582562 152688 582564 152697
rect 582616 152688 582618 152697
rect 582562 152623 582618 152632
rect 582562 149288 582618 149297
rect 582562 149223 582618 149232
rect 582576 149122 582604 149223
rect 582564 149116 582616 149122
rect 582564 149058 582616 149064
rect 2134 142216 2190 142225
rect 2134 142151 2190 142160
rect 2042 136776 2098 136785
rect 2042 136711 2098 136720
rect 110 126440 166 126449
rect 110 126375 166 126384
rect 124 111217 152 126375
rect 110 111208 166 111217
rect 110 111143 166 111152
rect 2042 110664 2098 110673
rect 2042 110599 2098 110608
rect 110 95024 166 95033
rect 110 94959 166 94968
rect 18 85232 74 85241
rect 18 85167 74 85176
rect 18 63608 74 63617
rect 18 63543 74 63552
rect 32 6769 60 63543
rect 124 59129 152 94959
rect 110 59120 166 59129
rect 110 59055 166 59064
rect 110 47832 166 47841
rect 110 47767 166 47776
rect 124 19961 152 47767
rect 2056 45529 2084 110599
rect 2148 97617 2176 142151
rect 582472 139392 582524 139398
rect 582470 139360 582472 139369
rect 582524 139360 582526 139369
rect 582470 139295 582526 139304
rect 582470 134600 582526 134609
rect 582470 134535 582526 134544
rect 582484 133958 582512 134535
rect 582472 133952 582524 133958
rect 582472 133894 582524 133900
rect 582380 126064 582432 126070
rect 582378 126032 582380 126041
rect 582432 126032 582434 126041
rect 582378 125967 582434 125976
rect 582378 119912 582434 119921
rect 582378 119847 582434 119856
rect 582392 118726 582420 119847
rect 582380 118720 582432 118726
rect 582380 118662 582432 118668
rect 582564 112872 582616 112878
rect 582562 112840 582564 112849
rect 582616 112840 582618 112849
rect 582562 112775 582618 112784
rect 582562 105360 582618 105369
rect 582562 105295 582618 105304
rect 582576 104922 582604 105295
rect 582564 104916 582616 104922
rect 582564 104858 582616 104864
rect 582472 99544 582524 99550
rect 582470 99512 582472 99521
rect 582524 99512 582526 99521
rect 582470 99447 582526 99456
rect 2134 97608 2190 97617
rect 2134 97543 2190 97552
rect 582470 90672 582526 90681
rect 582470 90607 582526 90616
rect 582484 89758 582512 90607
rect 582472 89752 582524 89758
rect 582472 89694 582524 89700
rect 582380 86216 582432 86222
rect 582378 86184 582380 86193
rect 582432 86184 582434 86193
rect 582378 86119 582434 86128
rect 2778 79248 2834 79257
rect 2778 79183 2834 79192
rect 2792 71641 2820 79183
rect 582378 76120 582434 76129
rect 582378 76055 582434 76064
rect 582392 75954 582420 76055
rect 582380 75948 582432 75954
rect 582380 75890 582432 75896
rect 582564 73024 582616 73030
rect 582562 72992 582564 73001
rect 582616 72992 582618 73001
rect 582562 72927 582618 72936
rect 2778 71632 2834 71641
rect 2778 71567 2834 71576
rect 582562 61432 582618 61441
rect 582562 61367 582618 61376
rect 582576 60790 582604 61367
rect 582564 60784 582616 60790
rect 582564 60726 582616 60732
rect 582472 59696 582524 59702
rect 582470 59664 582472 59673
rect 582524 59664 582526 59673
rect 582470 59599 582526 59608
rect 582654 46744 582710 46753
rect 582654 46679 582710 46688
rect 582380 46368 582432 46374
rect 582378 46336 582380 46345
rect 582432 46336 582434 46345
rect 582378 46271 582434 46280
rect 582668 46170 582696 46679
rect 582656 46164 582708 46170
rect 582656 46106 582708 46112
rect 2042 45520 2098 45529
rect 2042 45455 2098 45464
rect 582562 33144 582618 33153
rect 582562 33079 582564 33088
rect 582616 33079 582618 33088
rect 582564 33050 582616 33056
rect 582470 32192 582526 32201
rect 582470 32127 582526 32136
rect 582484 31822 582512 32127
rect 582472 31816 582524 31822
rect 582472 31758 582524 31764
rect 6056 29866 6084 30048
rect 11116 29866 11144 30048
rect 16176 29866 16204 30048
rect 21236 29866 21264 30048
rect 6012 29838 6084 29866
rect 11072 29838 11144 29866
rect 16132 29838 16204 29866
rect 21192 29838 21264 29866
rect 26296 29866 26324 30048
rect 31356 29866 31384 30048
rect 36416 29866 36444 30048
rect 41476 29866 41504 30048
rect 46536 29866 46564 30048
rect 51596 29866 51624 30048
rect 56656 29866 56684 30048
rect 61716 29866 61744 30048
rect 66776 29866 66804 30048
rect 71836 29866 71864 30048
rect 76896 29866 76924 30048
rect 81956 29866 81984 30048
rect 87016 29866 87044 30048
rect 92076 29866 92104 30048
rect 97136 29866 97164 30048
rect 102196 29866 102224 30048
rect 107256 29866 107284 30048
rect 112316 29866 112344 30048
rect 117376 29866 117404 30048
rect 122436 29866 122464 30048
rect 127496 29866 127524 30048
rect 132556 29866 132584 30048
rect 137616 29866 137644 30048
rect 142676 29866 142704 30048
rect 147736 29866 147764 30048
rect 152888 29866 152916 30048
rect 157948 29866 157976 30048
rect 163008 29866 163036 30048
rect 168068 29866 168096 30048
rect 173128 29866 173156 30048
rect 178188 29866 178216 30048
rect 183248 29866 183276 30048
rect 188308 29866 188336 30048
rect 193368 29866 193396 30048
rect 198428 29866 198456 30048
rect 203488 29866 203516 30048
rect 208548 29866 208576 30048
rect 213608 29866 213636 30048
rect 218668 29866 218696 30048
rect 223728 29866 223756 30048
rect 228788 29866 228816 30048
rect 233848 29866 233876 30048
rect 238908 29866 238936 30048
rect 243968 29866 243996 30048
rect 249028 29866 249056 30048
rect 254088 29866 254116 30048
rect 259148 29866 259176 30048
rect 264208 29866 264236 30048
rect 269268 29866 269296 30048
rect 274328 29866 274356 30048
rect 279388 29866 279416 30048
rect 284448 29866 284476 30048
rect 289508 29866 289536 30048
rect 294660 29866 294688 30048
rect 299720 29866 299748 30048
rect 26296 29838 26372 29866
rect 31356 29838 31432 29866
rect 36416 29838 36492 29866
rect 41476 29838 41552 29866
rect 46536 29838 46612 29866
rect 51596 29838 51672 29866
rect 56656 29838 56732 29866
rect 61716 29838 61792 29866
rect 66776 29838 66852 29866
rect 71836 29838 71912 29866
rect 76896 29838 76972 29866
rect 81956 29838 82032 29866
rect 6012 27606 6040 29838
rect 1308 27600 1360 27606
rect 1308 27542 1360 27548
rect 6000 27600 6052 27606
rect 6000 27542 6052 27548
rect 110 19952 166 19961
rect 110 19887 166 19896
rect 18 6760 74 6769
rect 18 6695 74 6704
rect 1320 3534 1348 27542
rect 11072 27062 11100 29838
rect 5448 27056 5500 27062
rect 5448 26998 5500 27004
rect 11060 27056 11112 27062
rect 11060 26998 11112 27004
rect 4068 26988 4120 26994
rect 4068 26930 4120 26936
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 584 480 612 3470
rect 1688 480 1716 4082
rect 2872 3460 2924 3466
rect 2872 3402 2924 3408
rect 2884 480 2912 3402
rect 4080 480 4108 26930
rect 5460 6914 5488 26998
rect 16132 26994 16160 29838
rect 16120 26988 16172 26994
rect 16120 26930 16172 26936
rect 21192 26926 21220 29838
rect 26344 27606 26372 29838
rect 26332 27600 26384 27606
rect 26332 27542 26384 27548
rect 29644 27600 29696 27606
rect 29644 27542 29696 27548
rect 6828 26920 6880 26926
rect 6828 26862 6880 26868
rect 21180 26920 21232 26926
rect 21180 26862 21232 26868
rect 6840 6914 6868 26862
rect 18604 25696 18656 25702
rect 18604 25638 18656 25644
rect 7564 25560 7616 25566
rect 7564 25502 7616 25508
rect 5276 6886 5488 6914
rect 6472 6886 6868 6914
rect 5276 480 5304 6886
rect 6472 480 6500 6886
rect 7576 4146 7604 25502
rect 11704 24132 11756 24138
rect 11704 24074 11756 24080
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7668 480 7696 4762
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8772 480 8800 3538
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 9956 2984 10008 2990
rect 9956 2926 10008 2932
rect 9968 480 9996 2926
rect 11164 480 11192 3470
rect 11716 2990 11744 24074
rect 14464 10328 14516 10334
rect 14464 10270 14516 10276
rect 12348 4888 12400 4894
rect 12348 4830 12400 4836
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 12360 480 12388 4830
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 13556 480 13584 3674
rect 14476 3466 14504 10270
rect 17040 6248 17092 6254
rect 17040 6190 17092 6196
rect 14738 3632 14794 3641
rect 14738 3567 14794 3576
rect 14464 3460 14516 3466
rect 14464 3402 14516 3408
rect 14752 480 14780 3567
rect 15934 3360 15990 3369
rect 15934 3295 15990 3304
rect 15948 480 15976 3295
rect 17052 480 17080 6190
rect 18616 3602 18644 25638
rect 29656 21418 29684 27542
rect 31404 27198 31432 29838
rect 36464 27606 36492 29838
rect 41524 27606 41552 29838
rect 46584 27606 46612 29838
rect 51644 27606 51672 29838
rect 56704 27606 56732 29838
rect 36452 27600 36504 27606
rect 36452 27542 36504 27548
rect 39304 27600 39356 27606
rect 39304 27542 39356 27548
rect 41512 27600 41564 27606
rect 41512 27542 41564 27548
rect 43444 27600 43496 27606
rect 43444 27542 43496 27548
rect 46572 27600 46624 27606
rect 46572 27542 46624 27548
rect 47584 27600 47636 27606
rect 47584 27542 47636 27548
rect 51632 27600 51684 27606
rect 51632 27542 51684 27548
rect 52368 27600 52420 27606
rect 52368 27542 52420 27548
rect 56692 27600 56744 27606
rect 56692 27542 56744 27548
rect 57888 27600 57940 27606
rect 57888 27542 57940 27548
rect 58624 27600 58676 27606
rect 58624 27542 58676 27548
rect 31392 27192 31444 27198
rect 31392 27134 31444 27140
rect 33784 27124 33836 27130
rect 33784 27066 33836 27072
rect 32404 27056 32456 27062
rect 32404 26998 32456 27004
rect 29644 21412 29696 21418
rect 29644 21354 29696 21360
rect 25504 19984 25556 19990
rect 25504 19926 25556 19932
rect 22744 13116 22796 13122
rect 22744 13058 22796 13064
rect 21824 6316 21876 6322
rect 21824 6258 21876 6264
rect 19432 3664 19484 3670
rect 19432 3606 19484 3612
rect 18604 3596 18656 3602
rect 18604 3538 18656 3544
rect 18236 3120 18288 3126
rect 18236 3062 18288 3068
rect 18248 480 18276 3062
rect 19444 480 19472 3606
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20640 480 20668 3538
rect 21836 480 21864 6258
rect 22756 3738 22784 13058
rect 23020 7948 23072 7954
rect 23020 7890 23072 7896
rect 22744 3732 22796 3738
rect 22744 3674 22796 3680
rect 23032 480 23060 7890
rect 24214 3768 24270 3777
rect 24214 3703 24270 3712
rect 24228 480 24256 3703
rect 25318 3496 25374 3505
rect 25318 3431 25374 3440
rect 25332 480 25360 3431
rect 25516 3126 25544 19926
rect 27712 9172 27764 9178
rect 27712 9114 27764 9120
rect 26516 6384 26568 6390
rect 26516 6326 26568 6332
rect 25504 3120 25556 3126
rect 25504 3062 25556 3068
rect 26528 480 26556 6326
rect 27724 480 27752 9114
rect 30104 6452 30156 6458
rect 30104 6394 30156 6400
rect 28908 3528 28960 3534
rect 28908 3470 28960 3476
rect 28920 480 28948 3470
rect 30116 480 30144 6394
rect 31300 3732 31352 3738
rect 31300 3674 31352 3680
rect 31312 480 31340 3674
rect 32416 3670 32444 26998
rect 33600 7812 33652 7818
rect 33600 7754 33652 7760
rect 32404 3664 32456 3670
rect 32404 3606 32456 3612
rect 32404 3256 32456 3262
rect 32404 3198 32456 3204
rect 32416 480 32444 3198
rect 33612 480 33640 7754
rect 33796 3534 33824 27066
rect 36544 26988 36596 26994
rect 36544 26930 36596 26936
rect 35164 26920 35216 26926
rect 35164 26862 35216 26868
rect 34796 3664 34848 3670
rect 34796 3606 34848 3612
rect 33784 3528 33836 3534
rect 33784 3470 33836 3476
rect 34808 480 34836 3606
rect 35176 3466 35204 26862
rect 36556 3602 36584 26930
rect 39316 11762 39344 27542
rect 40684 25764 40736 25770
rect 40684 25706 40736 25712
rect 39304 11756 39356 11762
rect 39304 11698 39356 11704
rect 39304 10396 39356 10402
rect 39304 10338 39356 10344
rect 37188 7880 37240 7886
rect 37188 7822 37240 7828
rect 36544 3596 36596 3602
rect 36544 3538 36596 3544
rect 35164 3460 35216 3466
rect 35164 3402 35216 3408
rect 35992 3392 36044 3398
rect 35992 3334 36044 3340
rect 36004 480 36032 3334
rect 37200 480 37228 7822
rect 39316 3670 39344 10338
rect 40696 3738 40724 25706
rect 41328 14476 41380 14482
rect 41328 14418 41380 14424
rect 40684 3732 40736 3738
rect 40684 3674 40736 3680
rect 39304 3664 39356 3670
rect 39304 3606 39356 3612
rect 39580 3596 39632 3602
rect 39580 3538 39632 3544
rect 38384 3324 38436 3330
rect 38384 3266 38436 3272
rect 38396 480 38424 3266
rect 39592 480 39620 3538
rect 41340 3534 41368 14418
rect 43168 7676 43220 7682
rect 43168 7618 43220 7624
rect 41880 3800 41932 3806
rect 41880 3742 41932 3748
rect 40684 3528 40736 3534
rect 40684 3470 40736 3476
rect 41328 3528 41380 3534
rect 41328 3470 41380 3476
rect 40696 480 40724 3470
rect 41892 480 41920 3742
rect 43076 3664 43128 3670
rect 43076 3606 43128 3612
rect 43088 480 43116 3606
rect 43180 3330 43208 7618
rect 43456 7614 43484 27542
rect 44272 9104 44324 9110
rect 44272 9046 44324 9052
rect 43444 7608 43496 7614
rect 43444 7550 43496 7556
rect 43168 3324 43220 3330
rect 43168 3266 43220 3272
rect 44284 480 44312 9046
rect 47596 6594 47624 27542
rect 50344 27192 50396 27198
rect 50344 27134 50396 27140
rect 49884 9036 49936 9042
rect 49884 8978 49936 8984
rect 47584 6588 47636 6594
rect 47584 6530 47636 6536
rect 47860 4956 47912 4962
rect 47860 4898 47912 4904
rect 45468 3868 45520 3874
rect 45468 3810 45520 3816
rect 45480 480 45508 3810
rect 46664 3732 46716 3738
rect 46664 3674 46716 3680
rect 46676 480 46704 3674
rect 47872 480 47900 4898
rect 48964 4208 49016 4214
rect 48964 4150 49016 4156
rect 48976 480 49004 4150
rect 49896 3874 49924 8978
rect 50160 8968 50212 8974
rect 50160 8910 50212 8916
rect 49884 3868 49936 3874
rect 49884 3810 49936 3816
rect 50172 480 50200 8910
rect 50356 7750 50384 27134
rect 52380 17270 52408 27542
rect 53104 27532 53156 27538
rect 53104 27474 53156 27480
rect 52368 17264 52420 17270
rect 52368 17206 52420 17212
rect 51724 15904 51776 15910
rect 51724 15846 51776 15852
rect 50344 7744 50396 7750
rect 50344 7686 50396 7692
rect 51356 5024 51408 5030
rect 51356 4966 51408 4972
rect 51368 480 51396 4966
rect 51736 3806 51764 15846
rect 52552 6180 52604 6186
rect 52552 6122 52604 6128
rect 51724 3800 51776 3806
rect 51724 3742 51776 3748
rect 52564 480 52592 6122
rect 53116 4214 53144 27474
rect 54484 25628 54536 25634
rect 54484 25570 54536 25576
rect 53104 4208 53156 4214
rect 53104 4150 53156 4156
rect 54496 3466 54524 25570
rect 57900 6526 57928 27542
rect 57888 6520 57940 6526
rect 57888 6462 57940 6468
rect 58440 5160 58492 5166
rect 58440 5102 58492 5108
rect 54944 5092 54996 5098
rect 54944 5034 54996 5040
rect 53748 3460 53800 3466
rect 53748 3402 53800 3408
rect 54484 3460 54536 3466
rect 54484 3402 54536 3408
rect 53760 480 53788 3402
rect 54956 480 54984 5034
rect 56048 4208 56100 4214
rect 56048 4150 56100 4156
rect 56060 480 56088 4150
rect 57244 3800 57296 3806
rect 57244 3742 57296 3748
rect 57256 480 57284 3742
rect 58452 480 58480 5102
rect 58636 4214 58664 27542
rect 61764 26234 61792 29838
rect 66824 27470 66852 29838
rect 66812 27464 66864 27470
rect 66812 27406 66864 27412
rect 69664 27464 69716 27470
rect 69664 27406 69716 27412
rect 68284 27396 68336 27402
rect 68284 27338 68336 27344
rect 65524 26852 65576 26858
rect 65524 26794 65576 26800
rect 61764 26206 62068 26234
rect 62040 18630 62068 26206
rect 62028 18624 62080 18630
rect 62028 18566 62080 18572
rect 63224 6656 63276 6662
rect 63224 6598 63276 6604
rect 62028 5228 62080 5234
rect 62028 5170 62080 5176
rect 59636 4412 59688 4418
rect 59636 4354 59688 4360
rect 58624 4208 58676 4214
rect 58624 4150 58676 4156
rect 59648 480 59676 4354
rect 60832 3868 60884 3874
rect 60832 3810 60884 3816
rect 60844 480 60872 3810
rect 62040 480 62068 5170
rect 63236 480 63264 6598
rect 65536 4418 65564 26794
rect 65616 5296 65668 5302
rect 65616 5238 65668 5244
rect 65524 4412 65576 4418
rect 65524 4354 65576 4360
rect 64328 3936 64380 3942
rect 64328 3878 64380 3884
rect 64340 480 64368 3878
rect 65628 2666 65656 5238
rect 68296 4214 68324 27338
rect 69676 15978 69704 27406
rect 71884 27334 71912 29838
rect 71872 27328 71924 27334
rect 71872 27270 71924 27276
rect 75184 27260 75236 27266
rect 75184 27202 75236 27208
rect 69664 15972 69716 15978
rect 69664 15914 69716 15920
rect 70308 11824 70360 11830
rect 70308 11766 70360 11772
rect 69112 5364 69164 5370
rect 69112 5306 69164 5312
rect 66720 4208 66772 4214
rect 66720 4150 66772 4156
rect 68284 4208 68336 4214
rect 68284 4150 68336 4156
rect 65536 2638 65656 2666
rect 65536 480 65564 2638
rect 66732 480 66760 4150
rect 67916 4004 67968 4010
rect 67916 3946 67968 3952
rect 67928 480 67956 3946
rect 69124 480 69152 5306
rect 70320 480 70348 11766
rect 72608 5432 72660 5438
rect 72608 5374 72660 5380
rect 71504 4072 71556 4078
rect 71504 4014 71556 4020
rect 71516 480 71544 4014
rect 72620 480 72648 5374
rect 75196 4758 75224 27202
rect 76944 26234 76972 29838
rect 82004 27470 82032 29838
rect 86972 29838 87044 29866
rect 92032 29838 92104 29866
rect 97092 29838 97164 29866
rect 102152 29838 102224 29866
rect 107212 29838 107284 29866
rect 112272 29838 112344 29866
rect 117332 29838 117404 29866
rect 122392 29838 122464 29866
rect 127452 29838 127524 29866
rect 132512 29838 132584 29866
rect 137572 29838 137644 29866
rect 142632 29838 142704 29866
rect 147692 29838 147764 29866
rect 152844 29838 152916 29866
rect 157904 29838 157976 29866
rect 162964 29838 163036 29866
rect 168024 29838 168096 29866
rect 173084 29838 173156 29866
rect 178144 29838 178216 29866
rect 183204 29838 183276 29866
rect 188264 29838 188336 29866
rect 193324 29838 193396 29866
rect 198384 29838 198456 29866
rect 203444 29838 203516 29866
rect 208504 29838 208576 29866
rect 213564 29838 213636 29866
rect 218624 29838 218696 29866
rect 223684 29838 223756 29866
rect 228744 29838 228816 29866
rect 233804 29838 233876 29866
rect 238864 29838 238936 29866
rect 243924 29838 243996 29866
rect 248984 29838 249056 29866
rect 254044 29838 254116 29866
rect 259104 29838 259176 29866
rect 264164 29838 264236 29866
rect 269224 29838 269296 29866
rect 274284 29838 274356 29866
rect 279344 29838 279416 29866
rect 284404 29838 284476 29866
rect 289464 29838 289536 29866
rect 294616 29838 294688 29866
rect 299676 29838 299748 29866
rect 304780 29850 304808 30048
rect 309840 29866 309868 30048
rect 314900 29866 314928 30048
rect 303620 29844 303672 29850
rect 81992 27464 82044 27470
rect 81992 27406 82044 27412
rect 83464 27464 83516 27470
rect 83464 27406 83516 27412
rect 82728 27192 82780 27198
rect 82728 27134 82780 27140
rect 79324 26784 79376 26790
rect 79324 26726 79376 26732
rect 76944 26206 77248 26234
rect 77220 6730 77248 26206
rect 77208 6724 77260 6730
rect 77208 6666 77260 6672
rect 76196 5500 76248 5506
rect 76196 5442 76248 5448
rect 73804 4752 73856 4758
rect 73804 4694 73856 4700
rect 75184 4752 75236 4758
rect 75184 4694 75236 4700
rect 73816 480 73844 4694
rect 75000 4140 75052 4146
rect 75000 4082 75052 4088
rect 75012 480 75040 4082
rect 76208 480 76236 5442
rect 79336 4214 79364 26726
rect 80888 6860 80940 6866
rect 80888 6802 80940 6808
rect 79692 4616 79744 4622
rect 79692 4558 79744 4564
rect 77392 4208 77444 4214
rect 77392 4150 77444 4156
rect 79324 4208 79376 4214
rect 79324 4150 79376 4156
rect 77404 480 77432 4150
rect 78588 3324 78640 3330
rect 78588 3266 78640 3272
rect 78600 480 78628 3266
rect 79704 480 79732 4558
rect 80900 480 80928 6802
rect 82740 3398 82768 27134
rect 83476 4758 83504 27406
rect 86776 27260 86828 27266
rect 86776 27202 86828 27208
rect 83464 4752 83516 4758
rect 83464 4694 83516 4700
rect 84476 4752 84528 4758
rect 84476 4694 84528 4700
rect 83280 4548 83332 4554
rect 83280 4490 83332 4496
rect 82084 3392 82136 3398
rect 82084 3334 82136 3340
rect 82728 3392 82780 3398
rect 82728 3334 82780 3340
rect 82096 480 82124 3334
rect 83292 480 83320 4490
rect 84488 480 84516 4694
rect 86788 3398 86816 27202
rect 86972 6866 87000 29838
rect 90364 27328 90416 27334
rect 90364 27270 90416 27276
rect 86960 6860 87012 6866
rect 86960 6802 87012 6808
rect 87972 6724 88024 6730
rect 87972 6666 88024 6672
rect 86868 4480 86920 4486
rect 86868 4422 86920 4428
rect 85672 3392 85724 3398
rect 85672 3334 85724 3340
rect 86776 3392 86828 3398
rect 86776 3334 86828 3340
rect 85684 480 85712 3334
rect 86880 480 86908 4422
rect 87984 480 88012 6666
rect 90376 4214 90404 27270
rect 92032 26790 92060 29838
rect 97092 27470 97120 29838
rect 102152 27470 102180 29838
rect 97080 27464 97132 27470
rect 97080 27406 97132 27412
rect 101404 27464 101456 27470
rect 101404 27406 101456 27412
rect 102140 27464 102192 27470
rect 102140 27406 102192 27412
rect 93768 27328 93820 27334
rect 93768 27270 93820 27276
rect 92020 26784 92072 26790
rect 92020 26726 92072 26732
rect 90456 4548 90508 4554
rect 90456 4490 90508 4496
rect 90364 4208 90416 4214
rect 90364 4150 90416 4156
rect 89168 3256 89220 3262
rect 89168 3198 89220 3204
rect 89180 480 89208 3198
rect 90468 2258 90496 4490
rect 91560 4208 91612 4214
rect 91560 4150 91612 4156
rect 90376 2230 90496 2258
rect 90376 480 90404 2230
rect 91572 480 91600 4150
rect 93780 3330 93808 27270
rect 98000 18624 98052 18630
rect 98000 18566 98052 18572
rect 98012 16574 98040 18566
rect 98012 16546 98224 16574
rect 94688 15972 94740 15978
rect 94688 15914 94740 15920
rect 93952 4480 94004 4486
rect 93952 4422 94004 4428
rect 92756 3324 92808 3330
rect 92756 3266 92808 3272
rect 93768 3324 93820 3330
rect 93768 3266 93820 3272
rect 92768 480 92796 3266
rect 93964 480 93992 4422
rect 94700 490 94728 15914
rect 97448 4412 97500 4418
rect 97448 4354 97500 4360
rect 96252 3188 96304 3194
rect 96252 3130 96304 3136
rect 94976 598 95188 626
rect 94976 490 95004 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 94700 462 95004 490
rect 95160 480 95188 598
rect 96264 480 96292 3130
rect 97460 480 97488 4354
rect 98196 490 98224 16546
rect 101416 11830 101444 27406
rect 107212 27402 107240 29838
rect 107200 27396 107252 27402
rect 107200 27338 107252 27344
rect 107568 27396 107620 27402
rect 107568 27338 107620 27344
rect 104900 17264 104952 17270
rect 104900 17206 104952 17212
rect 104912 16574 104940 17206
rect 104912 16546 105768 16574
rect 101404 11824 101456 11830
rect 101404 11766 101456 11772
rect 102232 6520 102284 6526
rect 102232 6462 102284 6468
rect 101036 4344 101088 4350
rect 101036 4286 101088 4292
rect 99840 3188 99892 3194
rect 99840 3130 99892 3136
rect 98472 598 98684 626
rect 98472 490 98500 598
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98196 462 98500 490
rect 98656 480 98684 598
rect 99852 480 99880 3130
rect 101048 480 101076 4286
rect 102244 480 102272 6462
rect 104532 4276 104584 4282
rect 104532 4218 104584 4224
rect 103336 3120 103388 3126
rect 103336 3062 103388 3068
rect 103348 480 103376 3062
rect 104544 480 104572 4218
rect 105740 480 105768 16546
rect 107580 3058 107608 27338
rect 112272 26234 112300 29838
rect 114468 27464 114520 27470
rect 114468 27406 114520 27412
rect 111812 26206 112300 26234
rect 111812 6662 111840 26206
rect 112812 7608 112864 7614
rect 112812 7550 112864 7556
rect 111800 6656 111852 6662
rect 111800 6598 111852 6604
rect 109316 6588 109368 6594
rect 109316 6530 109368 6536
rect 111616 6588 111668 6594
rect 111616 6530 111668 6536
rect 108120 6520 108172 6526
rect 108120 6462 108172 6468
rect 106924 3052 106976 3058
rect 106924 2994 106976 3000
rect 107568 3052 107620 3058
rect 107568 2994 107620 3000
rect 106936 480 106964 2994
rect 108132 480 108160 6462
rect 109328 480 109356 6530
rect 110512 3052 110564 3058
rect 110512 2994 110564 3000
rect 110524 480 110552 2994
rect 111628 480 111656 6530
rect 112824 480 112852 7550
rect 114480 2990 114508 27406
rect 117332 26858 117360 29838
rect 122392 27606 122420 29838
rect 127452 27606 127480 29838
rect 122380 27600 122432 27606
rect 122380 27542 122432 27548
rect 124864 27600 124916 27606
rect 124864 27542 124916 27548
rect 127440 27600 127492 27606
rect 127440 27542 127492 27548
rect 117320 26852 117372 26858
rect 117320 26794 117372 26800
rect 119988 22772 120040 22778
rect 119988 22714 120040 22720
rect 116400 11756 116452 11762
rect 116400 11698 116452 11704
rect 115204 6656 115256 6662
rect 115204 6598 115256 6604
rect 114008 2984 114060 2990
rect 114008 2926 114060 2932
rect 114468 2984 114520 2990
rect 114468 2926 114520 2932
rect 114020 480 114048 2926
rect 115216 480 115244 6598
rect 116412 480 116440 11698
rect 119896 7744 119948 7750
rect 119896 7686 119948 7692
rect 118792 2984 118844 2990
rect 118792 2926 118844 2932
rect 117596 2916 117648 2922
rect 117596 2858 117648 2864
rect 117608 480 117636 2858
rect 118804 480 118832 2926
rect 119908 480 119936 7686
rect 120000 2990 120028 22714
rect 122840 21412 122892 21418
rect 122840 21354 122892 21360
rect 122852 16574 122880 21354
rect 122852 16546 123064 16574
rect 122288 8016 122340 8022
rect 122288 7958 122340 7964
rect 119988 2984 120040 2990
rect 119988 2926 120040 2932
rect 121092 2916 121144 2922
rect 121092 2858 121144 2864
rect 121104 480 121132 2858
rect 122300 480 122328 7958
rect 123036 490 123064 16546
rect 124876 6186 124904 27542
rect 132512 27538 132540 29838
rect 132500 27532 132552 27538
rect 132500 27474 132552 27480
rect 137572 26234 137600 29838
rect 142632 26234 142660 29838
rect 136652 26206 137600 26234
rect 142172 26206 142660 26234
rect 125876 11756 125928 11762
rect 125876 11698 125928 11704
rect 124864 6180 124916 6186
rect 124864 6122 124916 6128
rect 124680 2848 124732 2854
rect 124680 2790 124732 2796
rect 123312 598 123524 626
rect 123312 490 123340 598
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123036 462 123340 490
rect 123496 480 123524 598
rect 124692 480 124720 2790
rect 125888 480 125916 11698
rect 136652 9042 136680 26206
rect 142172 15910 142200 26206
rect 142160 15904 142212 15910
rect 142160 15846 142212 15852
rect 144736 15904 144788 15910
rect 144736 15846 144788 15852
rect 136640 9036 136692 9042
rect 136640 8978 136692 8984
rect 141240 9036 141292 9042
rect 141240 8978 141292 8984
rect 132960 7744 133012 7750
rect 132960 7686 133012 7692
rect 129372 7608 129424 7614
rect 129372 7550 129424 7556
rect 129384 480 129412 7550
rect 132972 480 133000 7686
rect 136456 6180 136508 6186
rect 136456 6122 136508 6128
rect 136468 480 136496 6122
rect 141252 480 141280 8978
rect 144748 480 144776 15846
rect 147692 7682 147720 29838
rect 152844 26234 152872 29838
rect 157904 26234 157932 29838
rect 162964 27606 162992 29838
rect 168024 27606 168052 29838
rect 162124 27600 162176 27606
rect 162124 27542 162176 27548
rect 162952 27600 163004 27606
rect 162952 27542 163004 27548
rect 166264 27600 166316 27606
rect 166264 27542 166316 27548
rect 168012 27600 168064 27606
rect 168012 27542 168064 27548
rect 151832 26206 152872 26234
rect 157352 26206 157932 26234
rect 151832 10402 151860 26206
rect 157352 25770 157380 26206
rect 157340 25764 157392 25770
rect 157340 25706 157392 25712
rect 151820 10396 151872 10402
rect 151820 10338 151872 10344
rect 162136 9178 162164 27542
rect 162124 9172 162176 9178
rect 162124 9114 162176 9120
rect 166276 7954 166304 27542
rect 173084 26234 173112 29838
rect 178144 26234 178172 29838
rect 183204 26234 183232 29838
rect 188264 26234 188292 29838
rect 193324 27606 193352 29838
rect 190460 27600 190512 27606
rect 190460 27542 190512 27548
rect 193312 27600 193364 27606
rect 193312 27542 193364 27548
rect 172532 26206 173112 26234
rect 178052 26206 178172 26234
rect 182192 26206 183232 26234
rect 187712 26206 188292 26234
rect 172532 19990 172560 26206
rect 172520 19984 172572 19990
rect 172520 19926 172572 19932
rect 178052 13122 178080 26206
rect 182192 25702 182220 26206
rect 182180 25696 182232 25702
rect 182180 25638 182232 25644
rect 178040 13116 178092 13122
rect 178040 13058 178092 13064
rect 187712 8022 187740 26206
rect 190472 22778 190500 27542
rect 198384 26234 198412 29838
rect 203444 26234 203472 29838
rect 208504 26234 208532 29838
rect 213564 26234 213592 29838
rect 218624 26234 218652 29838
rect 223684 26234 223712 29838
rect 228744 26234 228772 29838
rect 233804 26234 233832 29838
rect 238864 26234 238892 29838
rect 243924 26234 243952 29838
rect 248984 26234 249012 29838
rect 254044 26234 254072 29838
rect 259104 26234 259132 29838
rect 264164 26234 264192 29838
rect 269224 26234 269252 29838
rect 274284 26234 274312 29838
rect 279344 26234 279372 29838
rect 284404 26234 284432 29838
rect 289464 26234 289492 29838
rect 294616 26234 294644 29838
rect 299676 26234 299704 29838
rect 303620 29786 303672 29792
rect 304768 29844 304820 29850
rect 304768 29786 304820 29792
rect 309796 29838 309868 29866
rect 314856 29838 314928 29866
rect 319960 29850 319988 30048
rect 325020 29866 325048 30048
rect 330080 29866 330108 30048
rect 318800 29844 318852 29850
rect 197372 26206 198412 26234
rect 202892 26206 203472 26234
rect 208412 26206 208532 26234
rect 212552 26206 213592 26234
rect 218072 26206 218652 26234
rect 223592 26206 223712 26234
rect 227732 26206 228772 26234
rect 233252 26206 233832 26234
rect 238772 26206 238892 26234
rect 242912 26206 243952 26234
rect 248432 26206 249012 26234
rect 253952 26206 254072 26234
rect 258092 26206 259132 26234
rect 263612 26206 264192 26234
rect 269132 26206 269252 26234
rect 273272 26206 274312 26234
rect 278792 26206 279372 26234
rect 284312 26206 284432 26234
rect 288452 26206 289492 26234
rect 293972 26206 294644 26234
rect 299492 26206 299704 26234
rect 190460 22772 190512 22778
rect 190460 22714 190512 22720
rect 187700 8016 187752 8022
rect 187700 7958 187752 7964
rect 166264 7948 166316 7954
rect 166264 7890 166316 7896
rect 147680 7676 147732 7682
rect 147680 7618 147732 7624
rect 148324 7676 148376 7682
rect 148324 7618 148376 7624
rect 148336 480 148364 7618
rect 197372 6662 197400 26206
rect 197360 6656 197412 6662
rect 197360 6598 197412 6604
rect 202892 6594 202920 26206
rect 202880 6588 202932 6594
rect 202880 6530 202932 6536
rect 208412 6526 208440 26206
rect 208400 6520 208452 6526
rect 208400 6462 208452 6468
rect 212552 4282 212580 26206
rect 218072 4350 218100 26206
rect 223592 4418 223620 26206
rect 227732 4486 227760 26206
rect 233252 4554 233280 26206
rect 238772 4622 238800 26206
rect 242912 4690 242940 26206
rect 248432 4758 248460 26206
rect 253952 5506 253980 26206
rect 253940 5500 253992 5506
rect 253940 5442 253992 5448
rect 258092 5438 258120 26206
rect 258080 5432 258132 5438
rect 258080 5374 258132 5380
rect 263612 5370 263640 26206
rect 263600 5364 263652 5370
rect 263600 5306 263652 5312
rect 269132 5302 269160 26206
rect 269120 5296 269172 5302
rect 269120 5238 269172 5244
rect 273272 5234 273300 26206
rect 273260 5228 273312 5234
rect 273260 5170 273312 5176
rect 278792 5166 278820 26206
rect 278780 5160 278832 5166
rect 278780 5102 278832 5108
rect 284312 5098 284340 26206
rect 284300 5092 284352 5098
rect 284300 5034 284352 5040
rect 288452 5030 288480 26206
rect 288440 5024 288492 5030
rect 288440 4966 288492 4972
rect 293972 4962 294000 26206
rect 299492 9110 299520 26206
rect 303632 14482 303660 29786
rect 309796 26234 309824 29838
rect 314856 27606 314884 29838
rect 318800 29786 318852 29792
rect 319948 29844 320000 29850
rect 319948 29786 320000 29792
rect 324976 29838 325048 29866
rect 330036 29838 330108 29866
rect 335140 29850 335168 30048
rect 333980 29844 334032 29850
rect 313924 27600 313976 27606
rect 313924 27542 313976 27548
rect 314844 27600 314896 27606
rect 314844 27542 314896 27548
rect 309152 26206 309824 26234
rect 303620 14476 303672 14482
rect 303620 14418 303672 14424
rect 299480 9104 299532 9110
rect 299480 9046 299532 9052
rect 309152 7886 309180 26206
rect 309140 7880 309192 7886
rect 309140 7822 309192 7828
rect 313936 7818 313964 27542
rect 313924 7812 313976 7818
rect 313924 7754 313976 7760
rect 318812 6458 318840 29786
rect 324976 26234 325004 29838
rect 330036 26234 330064 29838
rect 333980 29786 334032 29792
rect 335128 29844 335180 29850
rect 340200 29832 340228 30048
rect 345260 29866 345288 30048
rect 335128 29786 335180 29792
rect 340156 29804 340228 29832
rect 345216 29838 345288 29866
rect 350320 29850 350348 30048
rect 355380 29866 355408 30048
rect 360440 29866 360468 30048
rect 365500 29866 365528 30048
rect 370560 29866 370588 30048
rect 375620 29866 375648 30048
rect 349160 29844 349212 29850
rect 324332 26206 325004 26234
rect 329852 26206 330064 26234
rect 318800 6452 318852 6458
rect 318800 6394 318852 6400
rect 324332 6390 324360 26206
rect 324320 6384 324372 6390
rect 324320 6326 324372 6332
rect 329852 6322 329880 26206
rect 329840 6316 329892 6322
rect 329840 6258 329892 6264
rect 333992 6254 334020 29786
rect 340156 26234 340184 29804
rect 345216 26234 345244 29838
rect 349160 29786 349212 29792
rect 350308 29844 350360 29850
rect 350308 29786 350360 29792
rect 355336 29838 355408 29866
rect 360396 29838 360468 29866
rect 365456 29838 365528 29866
rect 370516 29838 370588 29866
rect 375576 29838 375648 29866
rect 380680 29850 380708 30048
rect 385740 29866 385768 30048
rect 390800 29866 390828 30048
rect 395860 29866 395888 30048
rect 400920 29866 400948 30048
rect 405980 29866 406008 30048
rect 411040 29866 411068 30048
rect 416100 29866 416128 30048
rect 421160 29866 421188 30048
rect 379520 29844 379572 29850
rect 339512 26206 340184 26234
rect 345032 26206 345244 26234
rect 333980 6248 334032 6254
rect 333980 6190 334032 6196
rect 293960 4956 294012 4962
rect 293960 4898 294012 4904
rect 339512 4894 339540 26206
rect 339500 4888 339552 4894
rect 339500 4830 339552 4836
rect 345032 4826 345060 26206
rect 345020 4820 345072 4826
rect 345020 4762 345072 4768
rect 248420 4752 248472 4758
rect 248420 4694 248472 4700
rect 242900 4684 242952 4690
rect 242900 4626 242952 4632
rect 238760 4616 238812 4622
rect 238760 4558 238812 4564
rect 233240 4548 233292 4554
rect 233240 4490 233292 4496
rect 227720 4480 227772 4486
rect 227720 4422 227772 4428
rect 223580 4412 223632 4418
rect 223580 4354 223632 4360
rect 218060 4344 218112 4350
rect 218060 4286 218112 4292
rect 212540 4276 212592 4282
rect 212540 4218 212592 4224
rect 349172 2854 349200 29786
rect 355336 26234 355364 29838
rect 360396 26234 360424 29838
rect 365456 27470 365484 29838
rect 365444 27464 365496 27470
rect 365444 27406 365496 27412
rect 370516 26234 370544 29838
rect 375576 27402 375604 29838
rect 379520 29786 379572 29792
rect 380668 29844 380720 29850
rect 380668 29786 380720 29792
rect 385696 29838 385768 29866
rect 390756 29838 390828 29866
rect 395816 29838 395888 29866
rect 400876 29838 400948 29866
rect 405936 29838 406008 29866
rect 410996 29838 411068 29866
rect 416056 29838 416128 29866
rect 421116 29838 421188 29866
rect 426220 29850 426248 30048
rect 431280 29866 431308 30048
rect 436432 29866 436460 30048
rect 425060 29844 425112 29850
rect 375564 27396 375616 27402
rect 375564 27338 375616 27344
rect 354692 26206 355364 26234
rect 360212 26206 360424 26234
rect 369872 26206 370544 26234
rect 354692 2922 354720 26206
rect 360212 2990 360240 26206
rect 369872 3058 369900 26206
rect 379532 3126 379560 29786
rect 385696 26234 385724 29838
rect 390756 26234 390784 29838
rect 395816 27334 395844 29838
rect 395804 27328 395856 27334
rect 395804 27270 395856 27276
rect 400876 26234 400904 29838
rect 405936 27266 405964 29838
rect 405924 27260 405976 27266
rect 405924 27202 405976 27208
rect 410996 27198 411024 29838
rect 410984 27192 411036 27198
rect 410984 27134 411036 27140
rect 416056 26234 416084 29838
rect 421116 26234 421144 29838
rect 425060 29786 425112 29792
rect 426208 29844 426260 29850
rect 426208 29786 426260 29792
rect 431236 29838 431308 29866
rect 436388 29838 436460 29866
rect 441492 29850 441520 30048
rect 440240 29844 440292 29850
rect 385052 26206 385724 26234
rect 390572 26206 390784 26234
rect 400232 26206 400904 26234
rect 415412 26206 416084 26234
rect 420932 26206 421144 26234
rect 385052 3194 385080 26206
rect 390572 3262 390600 26206
rect 400232 3330 400260 26206
rect 415412 3398 415440 26206
rect 420932 4146 420960 26206
rect 420920 4140 420972 4146
rect 420920 4082 420972 4088
rect 425072 4078 425100 29786
rect 431236 26234 431264 29838
rect 436388 26234 436416 29838
rect 440240 29786 440292 29792
rect 441480 29844 441532 29850
rect 446552 29832 446580 30048
rect 451612 29866 451640 30048
rect 456672 29866 456700 30048
rect 441480 29786 441532 29792
rect 446508 29804 446580 29832
rect 451568 29838 451640 29866
rect 456628 29838 456700 29866
rect 430592 26206 431264 26234
rect 436112 26206 436416 26234
rect 425060 4072 425112 4078
rect 425060 4014 425112 4020
rect 430592 4010 430620 26206
rect 430580 4004 430632 4010
rect 430580 3946 430632 3952
rect 436112 3942 436140 26206
rect 436100 3936 436152 3942
rect 436100 3878 436152 3884
rect 440252 3874 440280 29786
rect 446508 26234 446536 29804
rect 451568 26234 451596 29838
rect 456628 27606 456656 29838
rect 461732 29832 461760 30048
rect 466792 29832 466820 30048
rect 471852 29850 471880 30048
rect 476912 29866 476940 30048
rect 481972 29866 482000 30048
rect 487032 29866 487060 30048
rect 492092 29866 492120 30048
rect 497152 29866 497180 30048
rect 461688 29804 461760 29832
rect 466748 29804 466820 29832
rect 470600 29844 470652 29850
rect 454684 27600 454736 27606
rect 454684 27542 454736 27548
rect 456616 27600 456668 27606
rect 456616 27542 456668 27548
rect 445772 26206 446536 26234
rect 451292 26206 451596 26234
rect 440240 3868 440292 3874
rect 440240 3810 440292 3816
rect 445772 3806 445800 26206
rect 451292 25634 451320 26206
rect 451280 25628 451332 25634
rect 451280 25570 451332 25576
rect 454696 8974 454724 27542
rect 461688 26234 461716 29804
rect 466748 26234 466776 29804
rect 470600 29786 470652 29792
rect 471840 29844 471892 29850
rect 471840 29786 471892 29792
rect 476868 29838 476940 29866
rect 481928 29838 482000 29866
rect 486988 29838 487060 29866
rect 492048 29838 492120 29866
rect 497108 29838 497180 29866
rect 502212 29850 502240 30048
rect 507272 29866 507300 30048
rect 512332 29866 512360 30048
rect 517392 29866 517420 30048
rect 522452 29866 522480 30048
rect 527512 29866 527540 30048
rect 532572 29866 532600 30048
rect 537632 29866 537660 30048
rect 542692 29866 542720 30048
rect 500960 29844 501012 29850
rect 460952 26206 461716 26234
rect 466472 26206 466776 26234
rect 454684 8968 454736 8974
rect 454684 8910 454736 8916
rect 445760 3800 445812 3806
rect 445760 3742 445812 3748
rect 460952 3738 460980 26206
rect 460940 3732 460992 3738
rect 460940 3674 460992 3680
rect 466472 3670 466500 26206
rect 466460 3664 466512 3670
rect 466460 3606 466512 3612
rect 470612 3602 470640 29786
rect 476868 26234 476896 29838
rect 481928 26234 481956 29838
rect 486424 27192 486476 27198
rect 486424 27134 486476 27140
rect 476132 26206 476896 26234
rect 481652 26206 481956 26234
rect 470600 3596 470652 3602
rect 470600 3538 470652 3544
rect 476132 3534 476160 26206
rect 476120 3528 476172 3534
rect 476120 3470 476172 3476
rect 481652 3466 481680 26206
rect 486436 11762 486464 27134
rect 486988 27130 487016 29838
rect 486976 27124 487028 27130
rect 486976 27066 487028 27072
rect 492048 26234 492076 29838
rect 497108 27062 497136 29838
rect 500960 29786 501012 29792
rect 502200 29844 502252 29850
rect 502200 29786 502252 29792
rect 507228 29838 507300 29866
rect 512288 29838 512360 29866
rect 517348 29838 517420 29866
rect 522408 29838 522480 29866
rect 527468 29838 527540 29866
rect 532528 29838 532600 29866
rect 537588 29838 537660 29866
rect 542648 29838 542720 29866
rect 547752 29866 547780 30048
rect 552812 29866 552840 30048
rect 557872 29866 557900 30048
rect 547752 29838 547828 29866
rect 497096 27056 497148 27062
rect 497096 26998 497148 27004
rect 497464 27056 497516 27062
rect 497464 26998 497516 27004
rect 491312 26206 492076 26234
rect 486424 11756 486476 11762
rect 486424 11698 486476 11704
rect 491312 3777 491340 26206
rect 497476 7750 497504 26998
rect 497464 7744 497516 7750
rect 497464 7686 497516 7692
rect 491298 3768 491354 3777
rect 491298 3703 491354 3712
rect 500972 3641 501000 29786
rect 507228 26234 507256 29838
rect 512288 26234 512316 29838
rect 517348 27062 517376 29838
rect 517336 27056 517388 27062
rect 517336 26998 517388 27004
rect 518164 27056 518216 27062
rect 518164 26998 518216 27004
rect 506492 26206 507256 26234
rect 512012 26206 512316 26234
rect 506492 24138 506520 26206
rect 506480 24132 506532 24138
rect 506480 24074 506532 24080
rect 512012 6186 512040 26206
rect 518176 7682 518204 26998
rect 522408 26234 522436 29838
rect 527468 27130 527496 29838
rect 527456 27124 527508 27130
rect 527456 27066 527508 27072
rect 532528 27062 532556 29838
rect 532516 27056 532568 27062
rect 532516 26998 532568 27004
rect 537588 26234 537616 29838
rect 542648 26234 542676 29838
rect 521672 26206 522436 26234
rect 536852 26206 537616 26234
rect 542372 26206 542676 26234
rect 518164 7676 518216 7682
rect 518164 7618 518216 7624
rect 521672 7614 521700 26206
rect 536852 15910 536880 26206
rect 536840 15904 536892 15910
rect 536840 15846 536892 15852
rect 542372 9042 542400 26206
rect 542360 9036 542412 9042
rect 542360 8978 542412 8984
rect 521660 7608 521712 7614
rect 521660 7550 521712 7556
rect 512000 6180 512052 6186
rect 512000 6122 512052 6128
rect 500958 3632 501014 3641
rect 500958 3567 501014 3576
rect 547800 3466 547828 29838
rect 552768 29838 552840 29866
rect 557828 29838 557900 29866
rect 562932 29850 562960 30048
rect 567992 29866 568020 30048
rect 573052 29866 573080 30048
rect 578204 29866 578232 30048
rect 561680 29844 561732 29850
rect 552768 26234 552796 29838
rect 557828 26234 557856 29838
rect 561680 29786 561732 29792
rect 562920 29844 562972 29850
rect 562920 29786 562972 29792
rect 567948 29838 568020 29866
rect 573008 29838 573080 29866
rect 578160 29838 578232 29866
rect 552032 26206 552796 26234
rect 557552 26206 557856 26234
rect 552032 25566 552060 26206
rect 552020 25560 552072 25566
rect 552020 25502 552072 25508
rect 557552 10334 557580 26206
rect 557540 10328 557592 10334
rect 557540 10270 557592 10276
rect 561692 3505 561720 29786
rect 567948 26994 567976 29838
rect 567936 26988 567988 26994
rect 567936 26930 567988 26936
rect 573008 26234 573036 29838
rect 578160 26926 578188 29838
rect 578148 26920 578200 26926
rect 578148 26862 578200 26868
rect 572732 26206 573036 26234
rect 561678 3496 561734 3505
rect 481640 3460 481692 3466
rect 481640 3402 481692 3408
rect 547788 3460 547840 3466
rect 561678 3431 561734 3440
rect 547788 3402 547840 3408
rect 415400 3392 415452 3398
rect 572732 3369 572760 26206
rect 582656 19848 582708 19854
rect 582654 19816 582656 19825
rect 582708 19816 582710 19825
rect 582654 19751 582710 19760
rect 582472 6656 582524 6662
rect 582470 6624 582472 6633
rect 582524 6624 582526 6633
rect 582470 6559 582526 6568
rect 579804 3460 579856 3466
rect 579804 3402 579856 3408
rect 415400 3334 415452 3340
rect 572718 3360 572774 3369
rect 400220 3324 400272 3330
rect 572718 3295 572774 3304
rect 400220 3266 400272 3272
rect 390560 3256 390612 3262
rect 390560 3198 390612 3204
rect 385040 3188 385092 3194
rect 385040 3130 385092 3136
rect 379520 3120 379572 3126
rect 379520 3062 379572 3068
rect 369860 3052 369912 3058
rect 369860 2994 369912 3000
rect 360200 2984 360252 2990
rect 360200 2926 360252 2932
rect 354680 2916 354732 2922
rect 354680 2858 354732 2864
rect 349160 2848 349212 2854
rect 349160 2790 349212 2796
rect 579816 480 579844 3402
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 18 683712 74 683768
rect 582378 697196 582434 697232
rect 582378 697176 582380 697196
rect 582380 697176 582432 697196
rect 582432 697176 582434 697196
rect 582470 683868 582526 683904
rect 582470 683848 582472 683868
rect 582472 683848 582524 683868
rect 582524 683848 582526 683868
rect 110 676776 166 676832
rect 582378 676776 582434 676832
rect 2778 671200 2834 671256
rect 582378 670692 582380 670712
rect 582380 670692 582432 670712
rect 582432 670692 582434 670712
rect 582378 670656 582434 670692
rect 582470 662088 582526 662144
rect 2778 661136 2834 661192
rect 570 658180 572 658200
rect 572 658180 624 658200
rect 624 658180 626 658200
rect 570 658144 626 658180
rect 582378 647536 582434 647592
rect 18 645360 74 645416
rect 582378 644020 582434 644056
rect 582378 644000 582380 644020
rect 582380 644000 582432 644020
rect 582432 644000 582434 644020
rect 582378 632848 582434 632904
rect 570 632068 572 632088
rect 572 632068 624 632088
rect 624 632068 626 632088
rect 570 632032 626 632068
rect 582378 630828 582434 630864
rect 582378 630808 582380 630828
rect 582380 630808 582432 630828
rect 582432 630808 582434 630828
rect 110 629584 166 629640
rect 202 618568 258 618624
rect 582378 618196 582380 618216
rect 582380 618196 582432 618216
rect 582432 618196 582434 618216
rect 582378 618160 582434 618196
rect 582378 617500 582434 617536
rect 582378 617480 582380 617500
rect 582380 617480 582432 617500
rect 582432 617480 582434 617500
rect 202 613944 258 614000
rect 110 606600 166 606656
rect 582378 603608 582434 603664
rect 18 598168 74 598224
rect 580722 590960 580778 591016
rect 580722 588908 580778 588964
rect 110 582392 166 582448
rect 18 579672 74 579728
rect 582378 577652 582434 577688
rect 582378 577632 582380 577652
rect 582380 577632 582432 577652
rect 582432 577632 582434 577652
rect 582378 574232 582434 574288
rect 582378 564324 582434 564360
rect 582378 564304 582380 564324
rect 582380 564304 582432 564324
rect 582432 564304 582434 564324
rect 582378 559680 582434 559736
rect 110 554376 166 554432
rect 18 550976 74 551032
rect 582378 544856 582434 544912
rect 582378 537820 582380 537840
rect 582380 537820 582432 537840
rect 582432 537820 582434 537840
rect 582378 537784 582434 537820
rect 18 535200 74 535256
rect 582378 530168 582434 530224
rect 110 527312 166 527368
rect 582378 524492 582380 524512
rect 582380 524492 582432 524512
rect 582432 524492 582434 524512
rect 582378 524456 582434 524492
rect 2686 519424 2742 519480
rect 582378 515616 582434 515672
rect 2686 514800 2742 514856
rect 582378 511300 582380 511320
rect 582380 511300 582432 511320
rect 582432 511300 582434 511320
rect 582378 511264 582434 511300
rect 110 503920 166 503976
rect 18 502288 74 502344
rect 582378 500964 582380 500984
rect 582380 500964 582432 500984
rect 582432 500964 582434 500984
rect 582378 500928 582434 500964
rect 18 488144 74 488200
rect 582470 486240 582526 486296
rect 582378 484644 582380 484664
rect 582380 484644 582432 484664
rect 582432 484644 582434 484664
rect 582378 484608 582434 484644
rect 110 475088 166 475144
rect 2778 472368 2834 472424
rect 582562 471688 582618 471744
rect 582470 471452 582472 471472
rect 582472 471452 582524 471472
rect 582524 471452 582526 471472
rect 582470 471416 582526 471452
rect 2778 462576 2834 462632
rect 582562 458124 582564 458144
rect 582564 458124 582616 458144
rect 582616 458124 582618 458144
rect 582562 458088 582618 458124
rect 582378 457000 582434 457056
rect 110 456728 166 456784
rect 18 449792 74 449848
rect 582470 442312 582526 442368
rect 18 440952 74 441008
rect 582378 431604 582380 431624
rect 582380 431604 582432 431624
rect 582432 431604 582434 431624
rect 582378 431568 582434 431604
rect 582562 427760 582618 427816
rect 110 425176 166 425232
rect 2778 423544 2834 423600
rect 110 411032 166 411088
rect 582470 418276 582472 418296
rect 582472 418276 582524 418296
rect 582524 418276 582526 418296
rect 582470 418240 582526 418276
rect 582378 412936 582434 412992
rect 2778 409400 2834 409456
rect 582562 404948 582564 404968
rect 582564 404948 582616 404968
rect 582616 404948 582618 404968
rect 582562 404912 582618 404948
rect 582470 398384 582526 398440
rect 18 397976 74 398032
rect 110 393760 166 393816
rect 18 377984 74 378040
rect 18 358672 74 358728
rect 18 346568 74 346624
rect 582562 383716 582618 383752
rect 582562 383696 582564 383716
rect 582564 383696 582616 383716
rect 582616 383696 582618 383716
rect 582378 378428 582380 378448
rect 582380 378428 582432 378448
rect 582432 378428 582434 378448
rect 582378 378392 582434 378428
rect 2778 371320 2834 371376
rect 582378 369008 582434 369064
rect 582470 365100 582472 365120
rect 582472 365100 582524 365120
rect 582524 365100 582526 365120
rect 582470 365064 582526 365100
rect 2778 362208 2834 362264
rect 582654 354456 582710 354512
rect 582562 351908 582564 351928
rect 582564 351908 582616 351928
rect 582616 351908 582618 351928
rect 582562 351872 582618 351908
rect 110 345888 166 345944
rect 582562 339768 582618 339824
rect 110 330928 166 330984
rect 582378 325252 582380 325272
rect 582380 325252 582432 325272
rect 582432 325252 582434 325272
rect 582378 325216 582434 325252
rect 582470 325080 582526 325136
rect 2778 319232 2834 319288
rect 2778 315152 2834 315208
rect 582654 312060 582656 312080
rect 582656 312060 582708 312080
rect 582708 312060 582710 312080
rect 582654 312024 582710 312060
rect 582378 310548 582434 310584
rect 582378 310528 582380 310548
rect 582380 310528 582432 310548
rect 582432 310528 582434 310548
rect 110 306448 166 306504
rect 110 299376 166 299432
rect 18 293664 74 293720
rect 18 283600 74 283656
rect 18 254632 74 254688
rect 18 252184 74 252240
rect 582562 298732 582564 298752
rect 582564 298732 582616 298752
rect 582616 298732 582618 298752
rect 582562 298696 582618 298732
rect 582562 295840 582618 295896
rect 582654 281016 582710 281072
rect 582470 272212 582472 272232
rect 582472 272212 582524 272232
rect 582524 272212 582526 272232
rect 582470 272176 582526 272212
rect 582470 266464 582526 266520
rect 582378 258884 582380 258904
rect 582380 258884 582432 258904
rect 582432 258884 582434 258904
rect 582378 258848 582434 258884
rect 582378 251776 582434 251832
rect 582562 245556 582564 245576
rect 582564 245556 582616 245576
rect 582616 245556 582618 245576
rect 582562 245520 582618 245556
rect 110 241440 166 241496
rect 582746 237224 582802 237280
rect 110 236408 166 236464
rect 582654 232364 582656 232384
rect 582656 232364 582708 232384
rect 582708 232364 582710 232384
rect 582654 232328 582710 232364
rect 582654 222536 582710 222592
rect 2042 220768 2098 220824
rect 582470 219036 582472 219056
rect 582472 219036 582524 219056
rect 582524 219036 582526 219056
rect 582470 219000 582526 219036
rect 2042 214920 2098 214976
rect 582838 207848 582894 207904
rect 582378 205708 582380 205728
rect 582380 205708 582432 205728
rect 582432 205708 582434 205728
rect 582378 205672 582434 205708
rect 2042 204992 2098 205048
rect 110 202408 166 202464
rect 110 189352 166 189408
rect 18 189080 74 189136
rect 18 157936 74 157992
rect 110 150320 166 150376
rect 582562 193296 582618 193352
rect 582746 192516 582748 192536
rect 582748 192516 582800 192536
rect 582800 192516 582802 192536
rect 582746 192480 582802 192516
rect 582654 179188 582656 179208
rect 582656 179188 582708 179208
rect 582708 179188 582710 179208
rect 582654 179152 582710 179188
rect 582470 178608 582526 178664
rect 2778 173576 2834 173632
rect 582838 165860 582840 165880
rect 582840 165860 582892 165880
rect 582892 165860 582894 165880
rect 582838 165824 582894 165860
rect 582378 163920 582434 163976
rect 2778 162832 2834 162888
rect 582562 152668 582564 152688
rect 582564 152668 582616 152688
rect 582616 152668 582618 152688
rect 582562 152632 582618 152668
rect 582562 149232 582618 149288
rect 2134 142160 2190 142216
rect 2042 136720 2098 136776
rect 110 126384 166 126440
rect 110 111152 166 111208
rect 2042 110608 2098 110664
rect 110 94968 166 95024
rect 18 85176 74 85232
rect 18 63552 74 63608
rect 110 59064 166 59120
rect 110 47776 166 47832
rect 582470 139340 582472 139360
rect 582472 139340 582524 139360
rect 582524 139340 582526 139360
rect 582470 139304 582526 139340
rect 582470 134544 582526 134600
rect 582378 126012 582380 126032
rect 582380 126012 582432 126032
rect 582432 126012 582434 126032
rect 582378 125976 582434 126012
rect 582378 119856 582434 119912
rect 582562 112820 582564 112840
rect 582564 112820 582616 112840
rect 582616 112820 582618 112840
rect 582562 112784 582618 112820
rect 582562 105304 582618 105360
rect 582470 99492 582472 99512
rect 582472 99492 582524 99512
rect 582524 99492 582526 99512
rect 582470 99456 582526 99492
rect 2134 97552 2190 97608
rect 582470 90616 582526 90672
rect 582378 86164 582380 86184
rect 582380 86164 582432 86184
rect 582432 86164 582434 86184
rect 582378 86128 582434 86164
rect 2778 79192 2834 79248
rect 582378 76064 582434 76120
rect 582562 72972 582564 72992
rect 582564 72972 582616 72992
rect 582616 72972 582618 72992
rect 582562 72936 582618 72972
rect 2778 71576 2834 71632
rect 582562 61376 582618 61432
rect 582470 59644 582472 59664
rect 582472 59644 582524 59664
rect 582524 59644 582526 59664
rect 582470 59608 582526 59644
rect 582654 46688 582710 46744
rect 582378 46316 582380 46336
rect 582380 46316 582432 46336
rect 582432 46316 582434 46336
rect 582378 46280 582434 46316
rect 2042 45464 2098 45520
rect 582562 33108 582618 33144
rect 582562 33088 582564 33108
rect 582564 33088 582616 33108
rect 582616 33088 582618 33108
rect 582470 32136 582526 32192
rect 110 19896 166 19952
rect 18 6704 74 6760
rect 14738 3576 14794 3632
rect 15934 3304 15990 3360
rect 24214 3712 24270 3768
rect 25318 3440 25374 3496
rect 491298 3712 491354 3768
rect 500958 3576 501014 3632
rect 561678 3440 561734 3496
rect 582654 19796 582656 19816
rect 582656 19796 582708 19816
rect 582708 19796 582710 19816
rect 582654 19760 582710 19796
rect 582470 6604 582472 6624
rect 582472 6604 582524 6624
rect 582524 6604 582526 6624
rect 582470 6568 582526 6604
rect 572718 3304 572774 3360
<< metal3 >>
rect -960 697220 480 697460
rect 582373 697234 582439 697237
rect 583520 697234 584960 697324
rect 582373 697232 584960 697234
rect 582373 697176 582378 697232
rect 582434 697176 584960 697232
rect 582373 697174 584960 697176
rect 582373 697171 582439 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect -960 684254 674 684314
rect -960 684178 480 684254
rect 614 684178 674 684254
rect -960 684164 674 684178
rect 62 684118 674 684164
rect 62 683773 122 684118
rect 582465 683906 582531 683909
rect 583520 683906 584960 683996
rect 582465 683904 584960 683906
rect 582465 683848 582470 683904
rect 582526 683848 584960 683904
rect 582465 683846 584960 683848
rect 582465 683843 582531 683846
rect 13 683768 122 683773
rect 13 683712 18 683768
rect 74 683712 122 683768
rect 583520 683756 584960 683846
rect 13 683710 122 683712
rect 13 683707 79 683710
rect 105 676834 171 676837
rect 582373 676834 582439 676837
rect 105 676832 3434 676834
rect 105 676776 110 676832
rect 166 676806 3434 676832
rect 580766 676832 582439 676834
rect 580766 676806 582378 676832
rect 166 676776 4048 676806
rect 105 676774 4048 676776
rect 105 676771 171 676774
rect 3374 676746 4048 676774
rect 580244 676776 582378 676806
rect 582434 676776 582439 676832
rect 580244 676774 582439 676776
rect 580244 676746 580826 676774
rect 582373 676771 582439 676774
rect -960 671258 480 671348
rect 2773 671258 2839 671261
rect -960 671256 2839 671258
rect -960 671200 2778 671256
rect 2834 671200 2839 671256
rect -960 671198 2839 671200
rect -960 671108 480 671198
rect 2773 671195 2839 671198
rect 582373 670714 582439 670717
rect 583520 670714 584960 670804
rect 582373 670712 584960 670714
rect 582373 670656 582378 670712
rect 582434 670656 584960 670712
rect 582373 670654 584960 670656
rect 582373 670651 582439 670654
rect 583520 670564 584960 670654
rect 580244 662146 580826 662166
rect 582465 662146 582531 662149
rect 580244 662144 582531 662146
rect 580244 662106 582470 662144
rect 580766 662088 582470 662106
rect 582526 662088 582531 662144
rect 580766 662086 582531 662088
rect 582465 662083 582531 662086
rect 2773 661194 2839 661197
rect 2773 661192 3434 661194
rect 2773 661136 2778 661192
rect 2834 661190 3434 661192
rect 2834 661136 4048 661190
rect 2773 661134 4048 661136
rect 2773 661131 2839 661134
rect 3374 661130 4048 661134
rect -960 658202 480 658292
rect 565 658202 631 658205
rect -960 658200 631 658202
rect -960 658144 570 658200
rect 626 658144 631 658200
rect -960 658142 631 658144
rect -960 658052 480 658142
rect 565 658139 631 658142
rect 583520 657236 584960 657476
rect 582373 647594 582439 647597
rect 580766 647592 582439 647594
rect 580766 647536 582378 647592
rect 582434 647536 582439 647592
rect 580766 647534 582439 647536
rect 580766 647526 580826 647534
rect 582373 647531 582439 647534
rect 580244 647466 580826 647526
rect 13 645418 79 645421
rect 3374 645418 4048 645452
rect 13 645416 4048 645418
rect 13 645360 18 645416
rect 74 645392 4048 645416
rect 74 645360 3434 645392
rect 13 645358 3434 645360
rect 13 645355 79 645358
rect -960 644996 480 645236
rect 582373 644058 582439 644061
rect 583520 644058 584960 644148
rect 582373 644056 584960 644058
rect 582373 644000 582378 644056
rect 582434 644000 584960 644056
rect 582373 643998 584960 644000
rect 582373 643995 582439 643998
rect 583520 643908 584960 643998
rect 582373 632906 582439 632909
rect 580766 632904 582439 632906
rect 580766 632886 582378 632904
rect 580244 632848 582378 632886
rect 582434 632848 582439 632904
rect 580244 632846 582439 632848
rect 580244 632826 580826 632846
rect 582373 632843 582439 632846
rect -960 632090 480 632180
rect 565 632090 631 632093
rect -960 632088 631 632090
rect -960 632032 570 632088
rect 626 632032 631 632088
rect -960 632030 631 632032
rect -960 631940 480 632030
rect 565 632027 631 632030
rect 582373 630866 582439 630869
rect 583520 630866 584960 630956
rect 582373 630864 584960 630866
rect 582373 630808 582378 630864
rect 582434 630808 584960 630864
rect 582373 630806 584960 630808
rect 582373 630803 582439 630806
rect 583520 630716 584960 630806
rect 3742 629654 4048 629714
rect 105 629642 171 629645
rect 3742 629642 3802 629654
rect 105 629640 3802 629642
rect 105 629584 110 629640
rect 166 629584 3802 629640
rect 105 629582 3802 629584
rect 105 629579 171 629582
rect -960 619170 480 619260
rect -960 619110 674 619170
rect -960 619034 480 619110
rect 614 619034 674 619110
rect -960 619020 674 619034
rect 246 618974 674 619020
rect 246 618629 306 618974
rect 197 618624 306 618629
rect 197 618568 202 618624
rect 258 618568 306 618624
rect 197 618566 306 618568
rect 197 618563 263 618566
rect 580244 618218 580826 618246
rect 582373 618218 582439 618221
rect 580244 618216 582439 618218
rect 580244 618186 582378 618216
rect 580766 618160 582378 618186
rect 582434 618160 582439 618216
rect 580766 618158 582439 618160
rect 582373 618155 582439 618158
rect 582373 617538 582439 617541
rect 583520 617538 584960 617628
rect 582373 617536 584960 617538
rect 582373 617480 582378 617536
rect 582434 617480 584960 617536
rect 582373 617478 584960 617480
rect 582373 617475 582439 617478
rect 583520 617388 584960 617478
rect 197 614002 263 614005
rect 197 614000 3434 614002
rect 197 613944 202 614000
rect 258 613976 3434 614000
rect 258 613944 4048 613976
rect 197 613942 4048 613944
rect 197 613939 263 613942
rect 3374 613916 4048 613942
rect 105 606658 171 606661
rect 105 606656 306 606658
rect 105 606600 110 606656
rect 166 606600 306 606656
rect 105 606598 306 606600
rect 105 606595 171 606598
rect 246 606250 306 606598
rect 246 606204 674 606250
rect -960 606190 674 606204
rect -960 606114 480 606190
rect 614 606114 674 606190
rect -960 606054 674 606114
rect -960 605964 480 606054
rect 583520 604060 584960 604300
rect 582373 603666 582439 603669
rect 580766 603664 582439 603666
rect 580766 603608 582378 603664
rect 582434 603608 582439 603664
rect 580766 603606 582439 603608
rect 580244 603546 580826 603606
rect 582373 603603 582439 603606
rect 13 598226 79 598229
rect 3374 598226 4048 598238
rect 13 598224 4048 598226
rect 13 598168 18 598224
rect 74 598178 4048 598224
rect 74 598168 3434 598178
rect 13 598166 3434 598168
rect 13 598163 79 598166
rect -960 592908 480 593148
rect 580717 591018 580783 591021
rect 583520 591018 584960 591108
rect 580717 591016 584960 591018
rect 580717 590960 580722 591016
rect 580778 590960 584960 591016
rect 580717 590958 584960 590960
rect 580717 590955 580783 590958
rect 583520 590868 584960 590958
rect 580717 588966 580783 588969
rect 580244 588964 580783 588966
rect 580244 588908 580722 588964
rect 580778 588908 580783 588964
rect 580244 588906 580783 588908
rect 580717 588903 580783 588906
rect 105 582450 171 582453
rect 3374 582450 4048 582500
rect 105 582448 4048 582450
rect 105 582392 110 582448
rect 166 582440 4048 582448
rect 166 582392 3434 582440
rect 105 582390 3434 582392
rect 105 582387 171 582390
rect -960 580002 480 580092
rect -960 579942 674 580002
rect -960 579866 480 579942
rect 614 579866 674 579942
rect -960 579852 674 579866
rect 62 579806 674 579852
rect 62 579733 122 579806
rect 13 579728 122 579733
rect 13 579672 18 579728
rect 74 579672 122 579728
rect 13 579670 122 579672
rect 13 579667 79 579670
rect 582373 577690 582439 577693
rect 583520 577690 584960 577780
rect 582373 577688 584960 577690
rect 582373 577632 582378 577688
rect 582434 577632 584960 577688
rect 582373 577630 584960 577632
rect 582373 577627 582439 577630
rect 583520 577540 584960 577630
rect 580244 574290 580826 574326
rect 582373 574290 582439 574293
rect 580244 574288 582439 574290
rect 580244 574266 582378 574288
rect 580766 574232 582378 574266
rect 582434 574232 582439 574288
rect 580766 574230 582439 574232
rect 582373 574227 582439 574230
rect -960 566946 480 567036
rect -960 566886 3434 566946
rect -960 566796 480 566886
rect 3374 566762 3434 566886
rect 3374 566702 4048 566762
rect 582373 564362 582439 564365
rect 583520 564362 584960 564452
rect 582373 564360 584960 564362
rect 582373 564304 582378 564360
rect 582434 564304 584960 564360
rect 582373 564302 584960 564304
rect 582373 564299 582439 564302
rect 583520 564212 584960 564302
rect 582373 559738 582439 559741
rect 580766 559736 582439 559738
rect 580766 559686 582378 559736
rect 580244 559680 582378 559686
rect 582434 559680 582439 559736
rect 580244 559678 582439 559680
rect 580244 559626 580826 559678
rect 582373 559675 582439 559678
rect 105 554434 171 554437
rect 105 554432 306 554434
rect 105 554376 110 554432
rect 166 554376 306 554432
rect 105 554374 306 554376
rect 105 554371 171 554374
rect 246 554026 306 554374
rect 246 553980 674 554026
rect -960 553966 674 553980
rect -960 553890 480 553966
rect 614 553890 674 553966
rect -960 553830 674 553890
rect -960 553740 480 553830
rect 13 551034 79 551037
rect 13 551032 3434 551034
rect 13 550976 18 551032
rect 74 551024 3434 551032
rect 74 550976 4048 551024
rect 583520 551020 584960 551260
rect 13 550974 4048 550976
rect 13 550971 79 550974
rect 3374 550964 4048 550974
rect 580244 544914 580826 544924
rect 582373 544914 582439 544917
rect 580244 544912 582439 544914
rect 580244 544864 582378 544912
rect 580766 544856 582378 544864
rect 582434 544856 582439 544912
rect 580766 544854 582439 544856
rect 582373 544851 582439 544854
rect -960 540684 480 540924
rect 582373 537842 582439 537845
rect 583520 537842 584960 537932
rect 582373 537840 584960 537842
rect 582373 537784 582378 537840
rect 582434 537784 584960 537840
rect 582373 537782 584960 537784
rect 582373 537779 582439 537782
rect 583520 537692 584960 537782
rect 13 535258 79 535261
rect 3374 535258 4048 535286
rect 13 535256 4048 535258
rect 13 535200 18 535256
rect 74 535226 4048 535256
rect 74 535200 3434 535226
rect 13 535198 3434 535200
rect 13 535195 79 535198
rect 580244 530226 580826 530284
rect 582373 530226 582439 530229
rect 580244 530224 582439 530226
rect 580766 530168 582378 530224
rect 582434 530168 582439 530224
rect 580766 530166 582439 530168
rect 582373 530163 582439 530166
rect -960 527914 480 528004
rect -960 527854 674 527914
rect -960 527778 480 527854
rect 614 527778 674 527854
rect -960 527764 674 527778
rect 246 527718 674 527764
rect 105 527370 171 527373
rect 246 527370 306 527718
rect 105 527368 306 527370
rect 105 527312 110 527368
rect 166 527312 306 527368
rect 105 527310 306 527312
rect 105 527307 171 527310
rect 582373 524514 582439 524517
rect 583520 524514 584960 524604
rect 582373 524512 584960 524514
rect 582373 524456 582378 524512
rect 582434 524456 584960 524512
rect 582373 524454 584960 524456
rect 582373 524451 582439 524454
rect 583520 524364 584960 524454
rect 3742 519488 4048 519548
rect 2681 519482 2747 519485
rect 3742 519482 3802 519488
rect 2681 519480 3802 519482
rect 2681 519424 2686 519480
rect 2742 519424 3802 519480
rect 2681 519422 3802 519424
rect 2681 519419 2747 519422
rect 582373 515674 582439 515677
rect 580766 515672 582439 515674
rect 580766 515644 582378 515672
rect 580244 515616 582378 515644
rect 582434 515616 582439 515672
rect 580244 515614 582439 515616
rect 580244 515584 580826 515614
rect 582373 515611 582439 515614
rect -960 514858 480 514948
rect 2681 514858 2747 514861
rect -960 514856 2747 514858
rect -960 514800 2686 514856
rect 2742 514800 2747 514856
rect -960 514798 2747 514800
rect -960 514708 480 514798
rect 2681 514795 2747 514798
rect 582373 511322 582439 511325
rect 583520 511322 584960 511412
rect 582373 511320 584960 511322
rect 582373 511264 582378 511320
rect 582434 511264 584960 511320
rect 582373 511262 584960 511264
rect 582373 511259 582439 511262
rect 583520 511172 584960 511262
rect 105 503978 171 503981
rect 105 503976 3434 503978
rect 105 503920 110 503976
rect 166 503932 3434 503976
rect 166 503920 4048 503932
rect 105 503918 4048 503920
rect 105 503915 171 503918
rect 3374 503872 4048 503918
rect 13 502346 79 502349
rect 13 502344 122 502346
rect 13 502288 18 502344
rect 74 502288 122 502344
rect 13 502283 122 502288
rect 62 501938 122 502283
rect 62 501892 674 501938
rect -960 501878 674 501892
rect -960 501802 480 501878
rect 614 501802 674 501878
rect -960 501742 674 501802
rect -960 501652 480 501742
rect 580244 500986 580826 501004
rect 582373 500986 582439 500989
rect 580244 500984 582439 500986
rect 580244 500944 582378 500984
rect 580766 500928 582378 500944
rect 582434 500928 582439 500984
rect 580766 500926 582439 500928
rect 582373 500923 582439 500926
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 13 488202 79 488205
rect 13 488200 3434 488202
rect 13 488144 18 488200
rect 74 488194 3434 488200
rect 74 488144 4048 488194
rect 13 488142 4048 488144
rect 13 488139 79 488142
rect 3374 488134 4048 488142
rect 580244 486304 580826 486364
rect 580766 486298 580826 486304
rect 582465 486298 582531 486301
rect 580766 486296 582531 486298
rect 580766 486240 582470 486296
rect 582526 486240 582531 486296
rect 580766 486238 582531 486240
rect 582465 486235 582531 486238
rect 582373 484666 582439 484669
rect 583520 484666 584960 484756
rect 582373 484664 584960 484666
rect 582373 484608 582378 484664
rect 582434 484608 584960 484664
rect 582373 484606 584960 484608
rect 582373 484603 582439 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect -960 475630 674 475690
rect -960 475554 480 475630
rect 614 475554 674 475630
rect -960 475540 674 475554
rect 246 475494 674 475540
rect 105 475146 171 475149
rect 246 475146 306 475494
rect 105 475144 306 475146
rect 105 475088 110 475144
rect 166 475088 306 475144
rect 105 475086 306 475088
rect 105 475083 171 475086
rect 2773 472426 2839 472429
rect 3374 472426 4048 472456
rect 2773 472424 4048 472426
rect 2773 472368 2778 472424
rect 2834 472396 4048 472424
rect 2834 472368 3434 472396
rect 2773 472366 3434 472368
rect 2773 472363 2839 472366
rect 582557 471746 582623 471749
rect 580766 471744 582623 471746
rect 580766 471724 582562 471744
rect 580244 471688 582562 471724
rect 582618 471688 582623 471744
rect 580244 471686 582623 471688
rect 580244 471664 580826 471686
rect 582557 471683 582623 471686
rect 582465 471474 582531 471477
rect 583520 471474 584960 471564
rect 582465 471472 584960 471474
rect 582465 471416 582470 471472
rect 582526 471416 584960 471472
rect 582465 471414 584960 471416
rect 582465 471411 582531 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 2773 462634 2839 462637
rect -960 462632 2839 462634
rect -960 462576 2778 462632
rect 2834 462576 2839 462632
rect -960 462574 2839 462576
rect -960 462484 480 462574
rect 2773 462571 2839 462574
rect 582557 458146 582623 458149
rect 583520 458146 584960 458236
rect 582557 458144 584960 458146
rect 582557 458088 582562 458144
rect 582618 458088 584960 458144
rect 582557 458086 584960 458088
rect 582557 458083 582623 458086
rect 583520 457996 584960 458086
rect 580244 457058 580826 457084
rect 582373 457058 582439 457061
rect 580244 457056 582439 457058
rect 580244 457024 582378 457056
rect 580766 457000 582378 457024
rect 582434 457000 582439 457056
rect 580766 456998 582439 457000
rect 582373 456995 582439 456998
rect 105 456786 171 456789
rect 105 456784 3802 456786
rect 105 456728 110 456784
rect 166 456728 3802 456784
rect 105 456726 3802 456728
rect 105 456723 171 456726
rect 3742 456718 3802 456726
rect 3742 456658 4048 456718
rect 13 449850 79 449853
rect 13 449848 122 449850
rect 13 449792 18 449848
rect 74 449792 122 449848
rect 13 449787 122 449792
rect 62 449714 122 449787
rect 62 449668 674 449714
rect -960 449654 674 449668
rect -960 449578 480 449654
rect 614 449578 674 449654
rect -960 449518 674 449578
rect -960 449428 480 449518
rect 583520 444668 584960 444908
rect 580244 442384 580826 442444
rect 580766 442370 580826 442384
rect 582465 442370 582531 442373
rect 580766 442368 582531 442370
rect 580766 442312 582470 442368
rect 582526 442312 582531 442368
rect 580766 442310 582531 442312
rect 582465 442307 582531 442310
rect 13 441010 79 441013
rect 13 441008 3434 441010
rect 13 440952 18 441008
rect 74 440980 3434 441008
rect 74 440952 4048 440980
rect 13 440950 4048 440952
rect 13 440947 79 440950
rect 3374 440920 4048 440950
rect -960 436508 480 436748
rect 582373 431626 582439 431629
rect 583520 431626 584960 431716
rect 582373 431624 584960 431626
rect 582373 431568 582378 431624
rect 582434 431568 584960 431624
rect 582373 431566 584960 431568
rect 582373 431563 582439 431566
rect 583520 431476 584960 431566
rect 582557 427818 582623 427821
rect 580766 427816 582623 427818
rect 580766 427804 582562 427816
rect 580244 427760 582562 427804
rect 582618 427760 582623 427816
rect 580244 427758 582623 427760
rect 580244 427744 580826 427758
rect 582557 427755 582623 427758
rect 105 425234 171 425237
rect 3374 425234 4048 425242
rect 105 425232 4048 425234
rect 105 425176 110 425232
rect 166 425182 4048 425232
rect 166 425176 3434 425182
rect 105 425174 3434 425176
rect 105 425171 171 425174
rect -960 423602 480 423692
rect 2773 423602 2839 423605
rect -960 423600 2839 423602
rect -960 423544 2778 423600
rect 2834 423544 2839 423600
rect -960 423542 2839 423544
rect -960 423452 480 423542
rect 2773 423539 2839 423542
rect 582465 418298 582531 418301
rect 583520 418298 584960 418388
rect 582465 418296 584960 418298
rect 582465 418240 582470 418296
rect 582526 418240 584960 418296
rect 582465 418238 584960 418240
rect 582465 418235 582531 418238
rect 583520 418148 584960 418238
rect 580244 412994 580826 413042
rect 582373 412994 582439 412997
rect 580244 412992 582439 412994
rect 580244 412982 582378 412992
rect 580766 412936 582378 412982
rect 582434 412936 582439 412992
rect 580766 412934 582439 412936
rect 582373 412931 582439 412934
rect 105 411090 171 411093
rect 105 411088 306 411090
rect 105 411032 110 411088
rect 166 411032 306 411088
rect 105 411030 306 411032
rect 105 411027 171 411030
rect 246 410682 306 411030
rect 246 410636 674 410682
rect -960 410622 674 410636
rect -960 410546 480 410622
rect 614 410546 674 410622
rect -960 410486 674 410546
rect -960 410396 480 410486
rect 2773 409458 2839 409461
rect 3374 409458 4048 409504
rect 2773 409456 4048 409458
rect 2773 409400 2778 409456
rect 2834 409444 4048 409456
rect 2834 409400 3434 409444
rect 2773 409398 3434 409400
rect 2773 409395 2839 409398
rect 582557 404970 582623 404973
rect 583520 404970 584960 405060
rect 582557 404968 584960 404970
rect 582557 404912 582562 404968
rect 582618 404912 584960 404968
rect 582557 404910 584960 404912
rect 582557 404907 582623 404910
rect 583520 404820 584960 404910
rect 582465 398442 582531 398445
rect 580766 398440 582531 398442
rect 580766 398402 582470 398440
rect 580244 398384 582470 398402
rect 582526 398384 582531 398440
rect 580244 398382 582531 398384
rect 580244 398342 580826 398382
rect 582465 398379 582531 398382
rect 13 398034 79 398037
rect 13 398032 122 398034
rect 13 397976 18 398032
rect 74 397976 122 398032
rect 13 397971 122 397976
rect 62 397626 122 397971
rect 62 397580 674 397626
rect -960 397566 674 397580
rect -960 397490 480 397566
rect 614 397490 674 397566
rect -960 397430 674 397490
rect -960 397340 480 397430
rect 105 393818 171 393821
rect 105 393816 3434 393818
rect 105 393760 110 393816
rect 166 393766 3434 393816
rect 166 393760 4048 393766
rect 105 393758 4048 393760
rect 105 393755 171 393758
rect 3374 393706 4048 393758
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580244 383754 580826 383762
rect 582557 383754 582623 383757
rect 580244 383752 582623 383754
rect 580244 383702 582562 383752
rect 580766 383696 582562 383702
rect 582618 383696 582623 383752
rect 580766 383694 582623 383696
rect 582557 383691 582623 383694
rect 582373 378450 582439 378453
rect 583520 378450 584960 378540
rect 582373 378448 584960 378450
rect 582373 378392 582378 378448
rect 582434 378392 584960 378448
rect 582373 378390 584960 378392
rect 582373 378387 582439 378390
rect 583520 378300 584960 378390
rect 13 378042 79 378045
rect 13 378040 3434 378042
rect 13 377984 18 378040
rect 74 378028 3434 378040
rect 74 377984 4048 378028
rect 13 377982 4048 377984
rect 13 377979 79 377982
rect 3374 377968 4048 377982
rect -960 371378 480 371468
rect 2773 371378 2839 371381
rect -960 371376 2839 371378
rect -960 371320 2778 371376
rect 2834 371320 2839 371376
rect -960 371318 2839 371320
rect -960 371228 480 371318
rect 2773 371315 2839 371318
rect 580244 369066 580826 369122
rect 582373 369066 582439 369069
rect 580244 369064 582439 369066
rect 580244 369062 582378 369064
rect 580766 369008 582378 369062
rect 582434 369008 582439 369064
rect 580766 369006 582439 369008
rect 582373 369003 582439 369006
rect 582465 365122 582531 365125
rect 583520 365122 584960 365212
rect 582465 365120 584960 365122
rect 582465 365064 582470 365120
rect 582526 365064 584960 365120
rect 582465 365062 584960 365064
rect 582465 365059 582531 365062
rect 583520 364972 584960 365062
rect 2773 362266 2839 362269
rect 3374 362266 4048 362290
rect 2773 362264 4048 362266
rect 2773 362208 2778 362264
rect 2834 362230 4048 362264
rect 2834 362208 3434 362230
rect 2773 362206 3434 362208
rect 2773 362203 2839 362206
rect 13 358730 79 358733
rect 13 358728 122 358730
rect 13 358672 18 358728
rect 74 358672 122 358728
rect 13 358667 122 358672
rect 62 358594 122 358667
rect 62 358548 674 358594
rect -960 358534 674 358548
rect -960 358458 480 358534
rect 614 358458 674 358534
rect -960 358398 674 358458
rect -960 358308 480 358398
rect 582649 354514 582715 354517
rect 580766 354512 582715 354514
rect 580766 354482 582654 354512
rect 580244 354456 582654 354482
rect 582710 354456 582715 354512
rect 580244 354454 582715 354456
rect 580244 354422 580826 354454
rect 582649 354451 582715 354454
rect 582557 351930 582623 351933
rect 583520 351930 584960 352020
rect 582557 351928 584960 351930
rect 582557 351872 582562 351928
rect 582618 351872 584960 351928
rect 582557 351870 584960 351872
rect 582557 351867 582623 351870
rect 583520 351780 584960 351870
rect 13 346626 79 346629
rect 3374 346626 4048 346674
rect 13 346624 4048 346626
rect 13 346568 18 346624
rect 74 346614 4048 346624
rect 74 346568 3434 346614
rect 13 346566 3434 346568
rect 13 346563 79 346566
rect 105 345946 171 345949
rect 105 345944 306 345946
rect 105 345888 110 345944
rect 166 345888 306 345944
rect 105 345886 306 345888
rect 105 345883 171 345886
rect 246 345538 306 345886
rect 246 345492 674 345538
rect -960 345478 674 345492
rect -960 345402 480 345478
rect 614 345402 674 345478
rect -960 345342 674 345402
rect -960 345252 480 345342
rect 580244 339826 580826 339842
rect 582557 339826 582623 339829
rect 580244 339824 582623 339826
rect 580244 339782 582562 339824
rect 580766 339768 582562 339782
rect 582618 339768 582623 339824
rect 580766 339766 582623 339768
rect 582557 339763 582623 339766
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 105 330986 171 330989
rect 105 330984 3434 330986
rect 105 330928 110 330984
rect 166 330936 3434 330984
rect 166 330928 4048 330936
rect 105 330926 4048 330928
rect 105 330923 171 330926
rect 3374 330876 4048 330926
rect 582373 325274 582439 325277
rect 583520 325274 584960 325364
rect 582373 325272 584960 325274
rect 582373 325216 582378 325272
rect 582434 325216 584960 325272
rect 582373 325214 584960 325216
rect 582373 325211 582439 325214
rect 580244 325142 580826 325202
rect 580766 325138 580826 325142
rect 582465 325138 582531 325141
rect 580766 325136 582531 325138
rect 580766 325080 582470 325136
rect 582526 325080 582531 325136
rect 583520 325124 584960 325214
rect 580766 325078 582531 325080
rect 582465 325075 582531 325078
rect -960 319290 480 319380
rect 2773 319290 2839 319293
rect -960 319288 2839 319290
rect -960 319232 2778 319288
rect 2834 319232 2839 319288
rect -960 319230 2839 319232
rect -960 319140 480 319230
rect 2773 319227 2839 319230
rect 2773 315210 2839 315213
rect 2773 315208 3434 315210
rect 2773 315152 2778 315208
rect 2834 315198 3434 315208
rect 2834 315152 4048 315198
rect 2773 315150 4048 315152
rect 2773 315147 2839 315150
rect 3374 315138 4048 315150
rect 582649 312082 582715 312085
rect 583520 312082 584960 312172
rect 582649 312080 584960 312082
rect 582649 312024 582654 312080
rect 582710 312024 584960 312080
rect 582649 312022 584960 312024
rect 582649 312019 582715 312022
rect 583520 311932 584960 312022
rect 582373 310586 582439 310589
rect 580766 310584 582439 310586
rect 580766 310562 582378 310584
rect 580244 310528 582378 310562
rect 582434 310528 582439 310584
rect 580244 310526 582439 310528
rect 580244 310502 580826 310526
rect 582373 310523 582439 310526
rect 105 306506 171 306509
rect 62 306504 171 306506
rect 62 306448 110 306504
rect 166 306448 171 306504
rect 62 306443 171 306448
rect 62 306370 122 306443
rect 62 306324 674 306370
rect -960 306310 674 306324
rect -960 306234 480 306310
rect 614 306234 674 306310
rect -960 306174 674 306234
rect -960 306084 480 306174
rect 105 299434 171 299437
rect 3374 299434 4048 299460
rect 105 299432 4048 299434
rect 105 299376 110 299432
rect 166 299400 4048 299432
rect 166 299376 3434 299400
rect 105 299374 3434 299376
rect 105 299371 171 299374
rect 582557 298754 582623 298757
rect 583520 298754 584960 298844
rect 582557 298752 584960 298754
rect 582557 298696 582562 298752
rect 582618 298696 584960 298752
rect 582557 298694 584960 298696
rect 582557 298691 582623 298694
rect 583520 298604 584960 298694
rect 580244 295898 580826 295922
rect 582557 295898 582623 295901
rect 580244 295896 582623 295898
rect 580244 295862 582562 295896
rect 580766 295840 582562 295862
rect 582618 295840 582623 295896
rect 580766 295838 582623 295840
rect 582557 295835 582623 295838
rect 13 293722 79 293725
rect 13 293720 122 293722
rect 13 293664 18 293720
rect 74 293664 122 293720
rect 13 293659 122 293664
rect 62 293314 122 293659
rect 62 293268 674 293314
rect -960 293254 674 293268
rect -960 293178 480 293254
rect 614 293178 674 293254
rect -960 293118 674 293178
rect -960 293028 480 293118
rect 583520 285276 584960 285516
rect 3742 283662 4048 283722
rect 13 283658 79 283661
rect 3742 283658 3802 283662
rect 13 283656 3802 283658
rect 13 283600 18 283656
rect 74 283600 3802 283656
rect 13 283598 3802 283600
rect 13 283595 79 283598
rect 580244 281100 580826 281160
rect 580766 281074 580826 281100
rect 582649 281074 582715 281077
rect 580766 281072 582715 281074
rect 580766 281016 582654 281072
rect 582710 281016 582715 281072
rect 580766 281014 582715 281016
rect 582649 281011 582715 281014
rect -960 279972 480 280212
rect 582465 272234 582531 272237
rect 583520 272234 584960 272324
rect 582465 272232 584960 272234
rect 582465 272176 582470 272232
rect 582526 272176 584960 272232
rect 582465 272174 584960 272176
rect 582465 272171 582531 272174
rect 583520 272084 584960 272174
rect 3374 267924 4048 267984
rect 3374 267882 3434 267924
rect 430 267822 3434 267882
rect 430 267474 490 267822
rect 430 267414 674 267474
rect -960 267202 480 267292
rect 614 267202 674 267414
rect -960 267142 674 267202
rect -960 267052 480 267142
rect 582465 266522 582531 266525
rect 580766 266520 582531 266522
rect 580244 266464 582470 266520
rect 582526 266464 582531 266520
rect 580244 266462 582531 266464
rect 580244 266460 580826 266462
rect 582465 266459 582531 266462
rect 582373 258906 582439 258909
rect 583520 258906 584960 258996
rect 582373 258904 584960 258906
rect 582373 258848 582378 258904
rect 582434 258848 584960 258904
rect 582373 258846 584960 258848
rect 582373 258843 582439 258846
rect 583520 258756 584960 258846
rect 13 254690 79 254693
rect 13 254688 122 254690
rect 13 254632 18 254688
rect 74 254632 122 254688
rect 13 254627 122 254632
rect 62 254282 122 254627
rect 62 254236 674 254282
rect -960 254222 674 254236
rect -960 254146 480 254222
rect 614 254146 674 254222
rect -960 254086 674 254146
rect -960 253996 480 254086
rect 13 252242 79 252245
rect 3374 252242 4048 252246
rect 13 252240 4048 252242
rect 13 252184 18 252240
rect 74 252186 4048 252240
rect 74 252184 3434 252186
rect 13 252182 3434 252184
rect 13 252179 79 252182
rect 580244 251834 580826 251880
rect 582373 251834 582439 251837
rect 580244 251832 582439 251834
rect 580244 251820 582378 251832
rect 580766 251776 582378 251820
rect 582434 251776 582439 251832
rect 580766 251774 582439 251776
rect 582373 251771 582439 251774
rect 582557 245578 582623 245581
rect 583520 245578 584960 245668
rect 582557 245576 584960 245578
rect 582557 245520 582562 245576
rect 582618 245520 584960 245576
rect 582557 245518 584960 245520
rect 582557 245515 582623 245518
rect 583520 245428 584960 245518
rect 105 241498 171 241501
rect 105 241496 306 241498
rect 105 241440 110 241496
rect 166 241440 306 241496
rect 105 241438 306 241440
rect 105 241435 171 241438
rect 246 241226 306 241438
rect 246 241180 674 241226
rect -960 241166 674 241180
rect -960 241090 480 241166
rect 614 241090 674 241166
rect -960 241030 674 241090
rect -960 240940 480 241030
rect 582741 237282 582807 237285
rect 580766 237280 582807 237282
rect 580766 237240 582746 237280
rect 580244 237224 582746 237240
rect 582802 237224 582807 237280
rect 580244 237222 582807 237224
rect 580244 237180 580826 237222
rect 582741 237219 582807 237222
rect 105 236466 171 236469
rect 3374 236466 4048 236508
rect 105 236464 4048 236466
rect 105 236408 110 236464
rect 166 236448 4048 236464
rect 166 236408 3434 236448
rect 105 236406 3434 236408
rect 105 236403 171 236406
rect 582649 232386 582715 232389
rect 583520 232386 584960 232476
rect 582649 232384 584960 232386
rect 582649 232328 582654 232384
rect 582710 232328 584960 232384
rect 582649 232326 584960 232328
rect 582649 232323 582715 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580244 222594 580826 222600
rect 582649 222594 582715 222597
rect 580244 222592 582715 222594
rect 580244 222540 582654 222592
rect 580766 222536 582654 222540
rect 582710 222536 582715 222592
rect 580766 222534 582715 222536
rect 582649 222531 582715 222534
rect 2037 220826 2103 220829
rect 2037 220824 3434 220826
rect 2037 220768 2042 220824
rect 2098 220770 3434 220824
rect 2098 220768 4048 220770
rect 2037 220766 4048 220768
rect 2037 220763 2103 220766
rect 3374 220710 4048 220766
rect 582465 219058 582531 219061
rect 583520 219058 584960 219148
rect 582465 219056 584960 219058
rect 582465 219000 582470 219056
rect 582526 219000 584960 219056
rect 582465 218998 584960 219000
rect 582465 218995 582531 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 2037 214978 2103 214981
rect -960 214976 2103 214978
rect -960 214920 2042 214976
rect 2098 214920 2103 214976
rect -960 214918 2103 214920
rect -960 214828 480 214918
rect 2037 214915 2103 214918
rect 580244 207906 580826 207960
rect 582833 207906 582899 207909
rect 580244 207904 582899 207906
rect 580244 207900 582838 207904
rect 580766 207848 582838 207900
rect 582894 207848 582899 207904
rect 580766 207846 582899 207848
rect 582833 207843 582899 207846
rect 582373 205730 582439 205733
rect 583520 205730 584960 205820
rect 582373 205728 584960 205730
rect 582373 205672 582378 205728
rect 582434 205672 584960 205728
rect 582373 205670 584960 205672
rect 582373 205667 582439 205670
rect 583520 205580 584960 205670
rect 2037 205050 2103 205053
rect 2037 205048 3434 205050
rect 2037 204992 2042 205048
rect 2098 205032 3434 205048
rect 2098 204992 4048 205032
rect 2037 204990 4048 204992
rect 2037 204987 2103 204990
rect 3374 204972 4048 204990
rect 105 202466 171 202469
rect 105 202464 306 202466
rect 105 202408 110 202464
rect 166 202408 306 202464
rect 105 202406 306 202408
rect 105 202403 171 202406
rect 246 202058 306 202406
rect 246 202012 674 202058
rect -960 201998 674 202012
rect -960 201922 480 201998
rect 614 201922 674 201998
rect -960 201862 674 201922
rect -960 201772 480 201862
rect 582557 193354 582623 193357
rect 580766 193352 582623 193354
rect 580766 193320 582562 193352
rect 580244 193296 582562 193320
rect 582618 193296 582623 193352
rect 580244 193294 582623 193296
rect 580244 193260 580826 193294
rect 582557 193291 582623 193294
rect 582741 192538 582807 192541
rect 583520 192538 584960 192628
rect 582741 192536 584960 192538
rect 582741 192480 582746 192536
rect 582802 192480 584960 192536
rect 582741 192478 584960 192480
rect 582741 192475 582807 192478
rect 583520 192388 584960 192478
rect 105 189410 171 189413
rect 3374 189410 4048 189416
rect 105 189408 4048 189410
rect 105 189352 110 189408
rect 166 189356 4048 189408
rect 166 189352 3434 189356
rect 105 189350 3434 189352
rect 105 189347 171 189350
rect 13 189138 79 189141
rect 13 189136 122 189138
rect 13 189080 18 189136
rect 74 189080 122 189136
rect 13 189075 122 189080
rect 62 189002 122 189075
rect 62 188956 674 189002
rect -960 188942 674 188956
rect -960 188866 480 188942
rect 614 188866 674 188942
rect -960 188806 674 188866
rect -960 188716 480 188806
rect 582649 179210 582715 179213
rect 583520 179210 584960 179300
rect 582649 179208 584960 179210
rect 582649 179152 582654 179208
rect 582710 179152 584960 179208
rect 582649 179150 584960 179152
rect 582649 179147 582715 179150
rect 583520 179060 584960 179150
rect 580244 178666 580826 178680
rect 582465 178666 582531 178669
rect 580244 178664 582531 178666
rect 580244 178620 582470 178664
rect 580766 178608 582470 178620
rect 582526 178608 582531 178664
rect 580766 178606 582531 178608
rect 582465 178603 582531 178606
rect -960 175796 480 176036
rect 2773 173634 2839 173637
rect 3374 173634 4048 173678
rect 2773 173632 4048 173634
rect 2773 173576 2778 173632
rect 2834 173618 4048 173632
rect 2834 173576 3434 173618
rect 2773 173574 3434 173576
rect 2773 173571 2839 173574
rect 582833 165882 582899 165885
rect 583520 165882 584960 165972
rect 582833 165880 584960 165882
rect 582833 165824 582838 165880
rect 582894 165824 584960 165880
rect 582833 165822 584960 165824
rect 582833 165819 582899 165822
rect 583520 165732 584960 165822
rect 580244 163980 580826 164040
rect 580766 163978 580826 163980
rect 582373 163978 582439 163981
rect 580766 163976 582439 163978
rect 580766 163920 582378 163976
rect 582434 163920 582439 163976
rect 580766 163918 582439 163920
rect 582373 163915 582439 163918
rect -960 162890 480 162980
rect 2773 162890 2839 162893
rect -960 162888 2839 162890
rect -960 162832 2778 162888
rect 2834 162832 2839 162888
rect -960 162830 2839 162832
rect -960 162740 480 162830
rect 2773 162827 2839 162830
rect 13 157994 79 157997
rect 13 157992 3434 157994
rect 13 157936 18 157992
rect 74 157940 3434 157992
rect 74 157936 4048 157940
rect 13 157934 4048 157936
rect 13 157931 79 157934
rect 3374 157880 4048 157934
rect 582557 152690 582623 152693
rect 583520 152690 584960 152780
rect 582557 152688 584960 152690
rect 582557 152632 582562 152688
rect 582618 152632 584960 152688
rect 582557 152630 584960 152632
rect 582557 152627 582623 152630
rect 583520 152540 584960 152630
rect 105 150378 171 150381
rect 105 150376 306 150378
rect 105 150320 110 150376
rect 166 150320 306 150376
rect 105 150318 306 150320
rect 105 150315 171 150318
rect 246 149970 306 150318
rect 246 149924 674 149970
rect -960 149910 674 149924
rect -960 149834 480 149910
rect 614 149834 674 149910
rect -960 149774 674 149834
rect -960 149684 480 149774
rect 582557 149290 582623 149293
rect 580766 149288 582623 149290
rect 580766 149278 582562 149288
rect 580244 149232 582562 149278
rect 582618 149232 582623 149288
rect 580244 149230 582623 149232
rect 580244 149218 580826 149230
rect 582557 149227 582623 149230
rect 2129 142218 2195 142221
rect 2129 142216 3434 142218
rect 2129 142160 2134 142216
rect 2190 142202 3434 142216
rect 2190 142160 4048 142202
rect 2129 142158 4048 142160
rect 2129 142155 2195 142158
rect 3374 142142 4048 142158
rect 582465 139362 582531 139365
rect 583520 139362 584960 139452
rect 582465 139360 584960 139362
rect 582465 139304 582470 139360
rect 582526 139304 584960 139360
rect 582465 139302 584960 139304
rect 582465 139299 582531 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 2037 136778 2103 136781
rect -960 136776 2103 136778
rect -960 136720 2042 136776
rect 2098 136720 2103 136776
rect -960 136718 2103 136720
rect -960 136628 480 136718
rect 2037 136715 2103 136718
rect 580244 134602 580826 134638
rect 582465 134602 582531 134605
rect 580244 134600 582531 134602
rect 580244 134578 582470 134600
rect 580766 134544 582470 134578
rect 582526 134544 582531 134600
rect 580766 134542 582531 134544
rect 582465 134539 582531 134542
rect 105 126442 171 126445
rect 3374 126442 4048 126464
rect 105 126440 4048 126442
rect 105 126384 110 126440
rect 166 126404 4048 126440
rect 166 126384 3434 126404
rect 105 126382 3434 126384
rect 105 126379 171 126382
rect 582373 126034 582439 126037
rect 583520 126034 584960 126124
rect 582373 126032 584960 126034
rect 582373 125976 582378 126032
rect 582434 125976 584960 126032
rect 582373 125974 584960 125976
rect 582373 125971 582439 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 580244 119938 580826 119998
rect 580766 119914 580826 119938
rect 582373 119914 582439 119917
rect 580766 119912 582439 119914
rect 580766 119856 582378 119912
rect 582434 119856 582439 119912
rect 580766 119854 582439 119856
rect 582373 119851 582439 119854
rect 582557 112842 582623 112845
rect 583520 112842 584960 112932
rect 582557 112840 584960 112842
rect 582557 112784 582562 112840
rect 582618 112784 584960 112840
rect 582557 112782 584960 112784
rect 582557 112779 582623 112782
rect 583520 112692 584960 112782
rect 105 111210 171 111213
rect 105 111208 306 111210
rect 105 111152 110 111208
rect 166 111152 306 111208
rect 105 111150 306 111152
rect 105 111147 171 111150
rect 246 110802 306 111150
rect 246 110756 674 110802
rect -960 110742 674 110756
rect -960 110666 480 110742
rect 614 110666 674 110742
rect -960 110606 674 110666
rect 2037 110666 2103 110669
rect 3374 110666 4048 110726
rect 2037 110664 3434 110666
rect 2037 110608 2042 110664
rect 2098 110608 3434 110664
rect 2037 110606 3434 110608
rect -960 110516 480 110606
rect 2037 110603 2103 110606
rect 582557 105362 582623 105365
rect 580766 105360 582623 105362
rect 580766 105358 582562 105360
rect 580244 105304 582562 105358
rect 582618 105304 582623 105360
rect 580244 105302 582623 105304
rect 580244 105298 580826 105302
rect 582557 105299 582623 105302
rect 582465 99514 582531 99517
rect 583520 99514 584960 99604
rect 582465 99512 584960 99514
rect 582465 99456 582470 99512
rect 582526 99456 584960 99512
rect 582465 99454 584960 99456
rect 582465 99451 582531 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 2129 97610 2195 97613
rect -960 97608 2195 97610
rect -960 97552 2134 97608
rect 2190 97552 2195 97608
rect -960 97550 2195 97552
rect -960 97460 480 97550
rect 2129 97547 2195 97550
rect 105 95026 171 95029
rect 105 95024 3434 95026
rect 105 94968 110 95024
rect 166 94988 3434 95024
rect 166 94968 4048 94988
rect 105 94966 4048 94968
rect 105 94963 171 94966
rect 3374 94928 4048 94966
rect 580244 90674 580826 90718
rect 582465 90674 582531 90677
rect 580244 90672 582531 90674
rect 580244 90658 582470 90672
rect 580766 90616 582470 90658
rect 582526 90616 582531 90672
rect 580766 90614 582531 90616
rect 582465 90611 582531 90614
rect 582373 86186 582439 86189
rect 583520 86186 584960 86276
rect 582373 86184 584960 86186
rect 582373 86128 582378 86184
rect 582434 86128 584960 86184
rect 582373 86126 584960 86128
rect 582373 86123 582439 86126
rect 583520 86036 584960 86126
rect 13 85234 79 85237
rect 13 85232 122 85234
rect 13 85176 18 85232
rect 74 85176 122 85232
rect 13 85171 122 85176
rect 62 84826 122 85171
rect 62 84780 674 84826
rect -960 84766 674 84780
rect -960 84690 480 84766
rect 614 84690 674 84766
rect -960 84630 674 84690
rect -960 84540 480 84630
rect 2773 79250 2839 79253
rect 2773 79248 4048 79250
rect 2773 79192 2778 79248
rect 2834 79192 4048 79248
rect 2773 79190 4048 79192
rect 2773 79187 2839 79190
rect 582373 76122 582439 76125
rect 580766 76120 582439 76122
rect 580766 76078 582378 76120
rect 580244 76064 582378 76078
rect 582434 76064 582439 76120
rect 580244 76062 582439 76064
rect 580244 76018 580826 76062
rect 582373 76059 582439 76062
rect 582557 72994 582623 72997
rect 583520 72994 584960 73084
rect 582557 72992 584960 72994
rect 582557 72936 582562 72992
rect 582618 72936 584960 72992
rect 582557 72934 584960 72936
rect 582557 72931 582623 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 2773 71634 2839 71637
rect -960 71632 2839 71634
rect -960 71576 2778 71632
rect 2834 71576 2839 71632
rect -960 71574 2839 71576
rect -960 71484 480 71574
rect 2773 71571 2839 71574
rect 13 63610 79 63613
rect 13 63608 3802 63610
rect 13 63552 18 63608
rect 74 63552 3802 63608
rect 13 63550 3802 63552
rect 13 63547 79 63550
rect 3742 63512 3802 63550
rect 3742 63452 4048 63512
rect 580244 61434 580826 61438
rect 582557 61434 582623 61437
rect 580244 61432 582623 61434
rect 580244 61378 582562 61432
rect 580766 61376 582562 61378
rect 582618 61376 582623 61432
rect 580766 61374 582623 61376
rect 582557 61371 582623 61374
rect 582465 59666 582531 59669
rect 583520 59666 584960 59756
rect 582465 59664 584960 59666
rect 582465 59608 582470 59664
rect 582526 59608 584960 59664
rect 582465 59606 584960 59608
rect 582465 59603 582531 59606
rect 583520 59516 584960 59606
rect 105 59122 171 59125
rect 105 59120 306 59122
rect 105 59064 110 59120
rect 166 59064 306 59120
rect 105 59062 306 59064
rect 105 59059 171 59062
rect 246 58714 306 59062
rect 246 58668 674 58714
rect -960 58654 674 58668
rect -960 58578 480 58654
rect 614 58578 674 58654
rect -960 58518 674 58578
rect -960 58428 480 58518
rect 105 47834 171 47837
rect 105 47832 3434 47834
rect 105 47776 110 47832
rect 166 47776 3434 47832
rect 105 47774 3434 47776
rect 105 47771 171 47774
rect 3374 47714 4048 47774
rect 580244 46746 580826 46798
rect 582649 46746 582715 46749
rect 580244 46744 582715 46746
rect 580244 46738 582654 46744
rect 580766 46688 582654 46738
rect 582710 46688 582715 46744
rect 580766 46686 582715 46688
rect 582649 46683 582715 46686
rect 582373 46338 582439 46341
rect 583520 46338 584960 46428
rect 582373 46336 584960 46338
rect 582373 46280 582378 46336
rect 582434 46280 584960 46336
rect 582373 46278 584960 46280
rect 582373 46275 582439 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 2037 45522 2103 45525
rect -960 45520 2103 45522
rect -960 45464 2042 45520
rect 2098 45464 2103 45520
rect -960 45462 2103 45464
rect -960 45372 480 45462
rect 2037 45459 2103 45462
rect 582557 33146 582623 33149
rect 583520 33146 584960 33236
rect 582557 33144 584960 33146
rect 582557 33088 582562 33144
rect 582618 33088 584960 33144
rect 582557 33086 584960 33088
rect 582557 33083 582623 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect -960 32406 3434 32466
rect -960 32316 480 32406
rect 3374 32036 3434 32406
rect 582465 32194 582531 32197
rect 580766 32192 582531 32194
rect 580766 32158 582470 32192
rect 580244 32136 582470 32158
rect 582526 32136 582531 32192
rect 580244 32134 582531 32136
rect 580244 32098 580826 32134
rect 582465 32131 582531 32134
rect 3374 31976 4048 32036
rect 105 19954 171 19957
rect 105 19952 306 19954
rect 105 19896 110 19952
rect 166 19896 306 19952
rect 105 19894 306 19896
rect 105 19891 171 19894
rect 246 19546 306 19894
rect 582649 19818 582715 19821
rect 583520 19818 584960 19908
rect 582649 19816 584960 19818
rect 582649 19760 582654 19816
rect 582710 19760 584960 19816
rect 582649 19758 584960 19760
rect 582649 19755 582715 19758
rect 583520 19668 584960 19758
rect 246 19500 674 19546
rect -960 19486 674 19500
rect -960 19410 480 19486
rect 614 19410 674 19486
rect -960 19350 674 19410
rect -960 19260 480 19350
rect 13 6762 79 6765
rect 13 6760 122 6762
rect 13 6704 18 6760
rect 74 6704 122 6760
rect 13 6699 122 6704
rect 62 6626 122 6699
rect 582465 6626 582531 6629
rect 583520 6626 584960 6716
rect 62 6580 674 6626
rect -960 6566 674 6580
rect -960 6490 480 6566
rect 614 6490 674 6566
rect 582465 6624 584960 6626
rect 582465 6568 582470 6624
rect 582526 6568 584960 6624
rect 582465 6566 584960 6568
rect 582465 6563 582531 6566
rect -960 6430 674 6490
rect 583520 6476 584960 6566
rect -960 6340 480 6430
rect 24209 3770 24275 3773
rect 491293 3770 491359 3773
rect 24209 3768 491359 3770
rect 24209 3712 24214 3768
rect 24270 3712 491298 3768
rect 491354 3712 491359 3768
rect 24209 3710 491359 3712
rect 24209 3707 24275 3710
rect 491293 3707 491359 3710
rect 14733 3634 14799 3637
rect 500953 3634 501019 3637
rect 14733 3632 501019 3634
rect 14733 3576 14738 3632
rect 14794 3576 500958 3632
rect 501014 3576 501019 3632
rect 14733 3574 501019 3576
rect 14733 3571 14799 3574
rect 500953 3571 501019 3574
rect 25313 3498 25379 3501
rect 561673 3498 561739 3501
rect 25313 3496 561739 3498
rect 25313 3440 25318 3496
rect 25374 3440 561678 3496
rect 561734 3440 561739 3496
rect 25313 3438 561739 3440
rect 25313 3435 25379 3438
rect 561673 3435 561739 3438
rect 15929 3362 15995 3365
rect 572713 3362 572779 3365
rect 15929 3360 572779 3362
rect 15929 3304 15934 3360
rect 15990 3304 572718 3360
rect 572774 3304 572779 3360
rect 15929 3302 572779 3304
rect 15929 3299 15995 3302
rect 572713 3299 572779 3302
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 680788 2414 686898
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 680788 6134 690618
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 680788 9854 694338
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 680788 13574 698058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 680788 20414 705242
rect 23514 680788 24134 707162
rect 27234 680788 27854 709082
rect 30954 680788 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 680788 38414 686898
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 680788 42134 690618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 680788 45854 694338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 680788 49574 698058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 680788 56414 705242
rect 59514 680788 60134 707162
rect 63234 680788 63854 709082
rect 66954 680788 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 680788 74414 686898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 680788 78134 690618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 680788 81854 694338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 680788 85574 698058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 680788 92414 705242
rect 95514 680788 96134 707162
rect 99234 680788 99854 709082
rect 102954 680788 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 680788 110414 686898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 680788 114134 690618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 680788 117854 694338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 680788 121574 698058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 680788 128414 705242
rect 131514 680788 132134 707162
rect 135234 680788 135854 709082
rect 138954 680788 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 680788 146414 686898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 680788 150134 690618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 680788 153854 694338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 680788 157574 698058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 680788 164414 705242
rect 167514 680788 168134 707162
rect 171234 680788 171854 709082
rect 174954 680788 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 680788 182414 686898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 680788 186134 690618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 680788 189854 694338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 680788 193574 698058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 680788 200414 705242
rect 203514 680788 204134 707162
rect 207234 680788 207854 709082
rect 210954 680788 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 680788 218414 686898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 680788 222134 690618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 680788 225854 694338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 680788 229574 698058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 680788 236414 705242
rect 239514 680788 240134 707162
rect 243234 680788 243854 709082
rect 246954 680788 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 680788 254414 686898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 680788 258134 690618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 680788 261854 694338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 680788 265574 698058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 680788 272414 705242
rect 275514 680788 276134 707162
rect 279234 680788 279854 709082
rect 282954 680788 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 680788 290414 686898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 680788 294134 690618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 680788 297854 694338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 680788 301574 698058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 680788 308414 705242
rect 311514 680788 312134 707162
rect 315234 680788 315854 709082
rect 318954 680788 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 680788 326414 686898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 680788 330134 690618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 680788 333854 694338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 680788 337574 698058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 680788 344414 705242
rect 347514 680788 348134 707162
rect 351234 680788 351854 709082
rect 354954 680788 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 680788 362414 686898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 680788 366134 690618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 680788 369854 694338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 680788 373574 698058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 680788 380414 705242
rect 383514 680788 384134 707162
rect 387234 680788 387854 709082
rect 390954 680788 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 680788 398414 686898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 680788 402134 690618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 680788 405854 694338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 680788 409574 698058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 680788 416414 705242
rect 419514 680788 420134 707162
rect 423234 680788 423854 709082
rect 426954 680788 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 680788 434414 686898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 680788 438134 690618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 680788 441854 694338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 680788 445574 698058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 680788 452414 705242
rect 455514 680788 456134 707162
rect 459234 680788 459854 709082
rect 462954 680788 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 680788 470414 686898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 680788 474134 690618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 680788 477854 694338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 680788 481574 698058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 680788 488414 705242
rect 491514 680788 492134 707162
rect 495234 680788 495854 709082
rect 498954 680788 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 680788 506414 686898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 680788 510134 690618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 680788 513854 694338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 680788 517574 698058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 680788 524414 705242
rect 527514 680788 528134 707162
rect 531234 680788 531854 709082
rect 534954 680788 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 680788 542414 686898
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 680788 546134 690618
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 680788 549854 694338
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 680788 553574 698058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 680788 560414 705242
rect 563514 680788 564134 707162
rect 567234 680788 567854 709082
rect 570954 680788 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 680788 578414 686898
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 680788 582134 690618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 4400 669454 5000 669486
rect 4400 669218 4582 669454
rect 4818 669218 5000 669454
rect 4400 669134 5000 669218
rect 4400 668898 4582 669134
rect 4818 668898 5000 669134
rect 4400 668866 5000 668898
rect 127056 669454 127296 669486
rect 127056 669218 127058 669454
rect 127294 669218 127296 669454
rect 127056 669134 127296 669218
rect 127056 668898 127058 669134
rect 127294 668898 127296 669134
rect 127056 668866 127296 668898
rect 140294 669454 140534 669486
rect 140294 669218 140296 669454
rect 140532 669218 140534 669454
rect 140294 669134 140534 669218
rect 140294 668898 140296 669134
rect 140532 668898 140534 669134
rect 140294 668866 140534 668898
rect 147646 669454 147886 669486
rect 147646 669218 147648 669454
rect 147884 669218 147886 669454
rect 147646 669134 147886 669218
rect 147646 668898 147648 669134
rect 147884 668898 147886 669134
rect 147646 668866 147886 668898
rect 190318 669454 190558 669486
rect 190318 669218 190320 669454
rect 190556 669218 190558 669454
rect 190318 669134 190558 669218
rect 190318 668898 190320 669134
rect 190556 668898 190558 669134
rect 190318 668866 190558 668898
rect 229686 669454 229926 669486
rect 229686 669218 229688 669454
rect 229924 669218 229926 669454
rect 229686 669134 229926 669218
rect 229686 668898 229688 669134
rect 229924 668898 229926 669134
rect 229686 668866 229926 668898
rect 432438 669454 432678 669486
rect 432438 669218 432440 669454
rect 432676 669218 432678 669454
rect 432438 669134 432678 669218
rect 432438 668898 432440 669134
rect 432676 668898 432678 669134
rect 432438 668866 432678 668898
rect 439790 669454 440030 669486
rect 439790 669218 439792 669454
rect 440028 669218 440030 669454
rect 439790 669134 440030 669218
rect 439790 668898 439792 669134
rect 440028 668898 440030 669134
rect 439790 668866 440030 668898
rect 457008 669454 457248 669486
rect 457008 669218 457010 669454
rect 457246 669218 457248 669454
rect 457008 669134 457248 669218
rect 457008 668898 457010 669134
rect 457246 668898 457248 669134
rect 457008 668866 457248 668898
rect 579288 669454 579888 669486
rect 579288 669218 579470 669454
rect 579706 669218 579888 669454
rect 579288 669134 579888 669218
rect 579288 668898 579470 669134
rect 579706 668898 579888 669134
rect 579288 668866 579888 668898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect 5200 651454 5800 651486
rect 5200 651218 5382 651454
rect 5618 651218 5800 651454
rect 5200 651134 5800 651218
rect 5200 650898 5382 651134
rect 5618 650898 5800 651134
rect 5200 650866 5800 650898
rect 127456 651454 127696 651486
rect 127456 651218 127458 651454
rect 127694 651218 127696 651454
rect 127456 651134 127696 651218
rect 127456 650898 127458 651134
rect 127694 650898 127696 651134
rect 127456 650866 127696 650898
rect 140654 651454 140894 651486
rect 140654 651218 140656 651454
rect 140892 651218 140894 651454
rect 140654 651134 140894 651218
rect 140654 650898 140656 651134
rect 140892 650898 140894 651134
rect 140654 650866 140894 650898
rect 147286 651454 147526 651486
rect 147286 651218 147288 651454
rect 147524 651218 147526 651454
rect 147286 651134 147526 651218
rect 147286 650898 147288 651134
rect 147524 650898 147526 651134
rect 147286 650866 147526 650898
rect 149658 651454 149898 651486
rect 149658 651218 149660 651454
rect 149896 651218 149898 651454
rect 149658 651134 149898 651218
rect 149658 650898 149660 651134
rect 149896 650898 149898 651134
rect 149658 650866 149898 650898
rect 188306 651454 188546 651486
rect 188306 651218 188308 651454
rect 188544 651218 188546 651454
rect 188306 651134 188546 651218
rect 188306 650898 188308 651134
rect 188544 650898 188546 651134
rect 188306 650866 188546 650898
rect 190678 651454 190918 651486
rect 190678 651218 190680 651454
rect 190916 651218 190918 651454
rect 190678 651134 190918 651218
rect 190678 650898 190680 651134
rect 190916 650898 190918 651134
rect 190678 650866 190918 650898
rect 229326 651454 229566 651486
rect 229326 651218 229328 651454
rect 229564 651218 229566 651454
rect 229326 651134 229566 651218
rect 229326 650898 229328 651134
rect 229564 650898 229566 651134
rect 229326 650866 229566 650898
rect 230698 651454 230938 651486
rect 230698 651218 230700 651454
rect 230936 651218 230938 651454
rect 230698 651134 230938 651218
rect 230698 650898 230700 651134
rect 230936 650898 230938 651134
rect 230698 650866 230938 650898
rect 269346 651454 269586 651486
rect 269346 651218 269348 651454
rect 269584 651218 269586 651454
rect 269346 651134 269586 651218
rect 269346 650898 269348 651134
rect 269584 650898 269586 651134
rect 269346 650866 269586 650898
rect 270718 651454 270958 651486
rect 270718 651218 270720 651454
rect 270956 651218 270958 651454
rect 270718 651134 270958 651218
rect 270718 650898 270720 651134
rect 270956 650898 270958 651134
rect 270718 650866 270958 650898
rect 309366 651454 309606 651486
rect 309366 651218 309368 651454
rect 309604 651218 309606 651454
rect 309366 651134 309606 651218
rect 309366 650898 309368 651134
rect 309604 650898 309606 651134
rect 309366 650866 309606 650898
rect 310562 651454 310802 651486
rect 310562 651218 310564 651454
rect 310800 651218 310802 651454
rect 310562 651134 310802 651218
rect 310562 650898 310564 651134
rect 310800 650898 310802 651134
rect 310562 650866 310802 650898
rect 311738 651454 311978 651486
rect 311738 651218 311740 651454
rect 311976 651218 311978 651454
rect 311738 651134 311978 651218
rect 311738 650898 311740 651134
rect 311976 650898 311978 651134
rect 311738 650866 311978 650898
rect 350386 651454 350626 651486
rect 350386 651218 350388 651454
rect 350624 651218 350626 651454
rect 350386 651134 350626 651218
rect 350386 650898 350388 651134
rect 350624 650898 350626 651134
rect 350386 650866 350626 650898
rect 352758 651454 352998 651486
rect 352758 651218 352760 651454
rect 352996 651218 352998 651454
rect 352758 651134 352998 651218
rect 352758 650898 352760 651134
rect 352996 650898 352998 651134
rect 352758 650866 352998 650898
rect 391406 651454 391646 651486
rect 391406 651218 391408 651454
rect 391644 651218 391646 651454
rect 391406 651134 391646 651218
rect 391406 650898 391408 651134
rect 391644 650898 391646 651134
rect 391406 650866 391646 650898
rect 392778 651454 393018 651486
rect 392778 651218 392780 651454
rect 393016 651218 393018 651454
rect 392778 651134 393018 651218
rect 392778 650898 392780 651134
rect 393016 650898 393018 651134
rect 392778 650866 393018 650898
rect 431426 651454 431666 651486
rect 431426 651218 431428 651454
rect 431664 651218 431666 651454
rect 431426 651134 431666 651218
rect 431426 650898 431428 651134
rect 431664 650898 431666 651134
rect 431426 650866 431666 650898
rect 432798 651454 433038 651486
rect 432798 651218 432800 651454
rect 433036 651218 433038 651454
rect 432798 651134 433038 651218
rect 432798 650898 432800 651134
rect 433036 650898 433038 651134
rect 432798 650866 433038 650898
rect 439430 651454 439670 651486
rect 439430 651218 439432 651454
rect 439668 651218 439670 651454
rect 439430 651134 439670 651218
rect 439430 650898 439432 651134
rect 439668 650898 439670 651134
rect 439430 650866 439670 650898
rect 456608 651454 456848 651486
rect 456608 651218 456610 651454
rect 456846 651218 456848 651454
rect 456608 651134 456848 651218
rect 456608 650898 456610 651134
rect 456846 650898 456848 651134
rect 456608 650866 456848 650898
rect 578488 651454 579088 651486
rect 578488 651218 578670 651454
rect 578906 651218 579088 651454
rect 578488 651134 579088 651218
rect 578488 650898 578670 651134
rect 578906 650898 579088 651134
rect 578488 650866 579088 650898
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 4400 633454 5000 633486
rect 4400 633218 4582 633454
rect 4818 633218 5000 633454
rect 4400 633134 5000 633218
rect 4400 632898 4582 633134
rect 4818 632898 5000 633134
rect 4400 632866 5000 632898
rect 12296 633454 12644 633486
rect 12296 633218 12352 633454
rect 12588 633218 12644 633454
rect 12296 633134 12644 633218
rect 12296 632898 12352 633134
rect 12588 632898 12644 633134
rect 12296 632866 12644 632898
rect 107360 633454 107708 633486
rect 107360 633218 107416 633454
rect 107652 633218 107708 633454
rect 107360 633134 107708 633218
rect 107360 632898 107416 633134
rect 107652 632898 107708 633134
rect 107360 632866 107708 632898
rect 127056 633454 127296 633486
rect 127056 633218 127058 633454
rect 127294 633218 127296 633454
rect 127056 633134 127296 633218
rect 127056 632898 127058 633134
rect 127294 632898 127296 633134
rect 127056 632866 127296 632898
rect 140294 633454 140534 633486
rect 140294 633218 140296 633454
rect 140532 633218 140534 633454
rect 140294 633134 140534 633218
rect 140294 632898 140296 633134
rect 140532 632898 140534 633134
rect 140294 632866 140534 632898
rect 141100 633454 141340 633486
rect 141100 633218 141102 633454
rect 141338 633218 141340 633454
rect 141100 633134 141340 633218
rect 141100 632898 141102 633134
rect 141338 632898 141340 633134
rect 141100 632866 141340 632898
rect 147646 633454 147886 633486
rect 147646 633218 147648 633454
rect 147884 633218 147886 633454
rect 147646 633134 147886 633218
rect 147646 632898 147648 633134
rect 147884 632898 147886 633134
rect 147646 632866 147886 632898
rect 149298 633454 149538 633486
rect 149298 633218 149300 633454
rect 149536 633218 149538 633454
rect 149298 633134 149538 633218
rect 149298 632898 149300 633134
rect 149536 632898 149538 633134
rect 149298 632866 149538 632898
rect 150104 633454 150344 633486
rect 150104 633218 150106 633454
rect 150342 633218 150344 633454
rect 150104 633134 150344 633218
rect 150104 632898 150106 633134
rect 150342 632898 150344 633134
rect 150104 632866 150344 632898
rect 159104 633454 159344 633486
rect 159104 633218 159106 633454
rect 159342 633218 159344 633454
rect 159104 633134 159344 633218
rect 159104 632898 159106 633134
rect 159342 632898 159344 633134
rect 159104 632866 159344 632898
rect 168104 633454 168344 633486
rect 168104 633218 168106 633454
rect 168342 633218 168344 633454
rect 168104 633134 168344 633218
rect 168104 632898 168106 633134
rect 168342 632898 168344 633134
rect 168104 632866 168344 632898
rect 177104 633454 177344 633486
rect 177104 633218 177106 633454
rect 177342 633218 177344 633454
rect 177104 633134 177344 633218
rect 177104 632898 177106 633134
rect 177342 632898 177344 633134
rect 177104 632866 177344 632898
rect 186104 633454 186344 633486
rect 186104 633218 186106 633454
rect 186342 633218 186344 633454
rect 186104 633134 186344 633218
rect 186104 632898 186106 633134
rect 186342 632898 186344 633134
rect 186104 632866 186344 632898
rect 188666 633454 188906 633486
rect 188666 633218 188668 633454
rect 188904 633218 188906 633454
rect 188666 633134 188906 633218
rect 188666 632898 188668 633134
rect 188904 632898 188906 633134
rect 188666 632866 188906 632898
rect 190318 633454 190558 633486
rect 190318 633218 190320 633454
rect 190556 633218 190558 633454
rect 190318 633134 190558 633218
rect 190318 632898 190320 633134
rect 190556 632898 190558 633134
rect 190318 632866 190558 632898
rect 191124 633454 191364 633486
rect 191124 633218 191126 633454
rect 191362 633218 191364 633454
rect 191124 633134 191364 633218
rect 191124 632898 191126 633134
rect 191362 632898 191364 633134
rect 191124 632866 191364 632898
rect 200124 633454 200364 633486
rect 200124 633218 200126 633454
rect 200362 633218 200364 633454
rect 200124 633134 200364 633218
rect 200124 632898 200126 633134
rect 200362 632898 200364 633134
rect 200124 632866 200364 632898
rect 209124 633454 209364 633486
rect 209124 633218 209126 633454
rect 209362 633218 209364 633454
rect 209124 633134 209364 633218
rect 209124 632898 209126 633134
rect 209362 632898 209364 633134
rect 209124 632866 209364 632898
rect 218124 633454 218364 633486
rect 218124 633218 218126 633454
rect 218362 633218 218364 633454
rect 218124 633134 218364 633218
rect 218124 632898 218126 633134
rect 218362 632898 218364 633134
rect 218124 632866 218364 632898
rect 227124 633454 227364 633486
rect 227124 633218 227126 633454
rect 227362 633218 227364 633454
rect 227124 633134 227364 633218
rect 227124 632898 227126 633134
rect 227362 632898 227364 633134
rect 227124 632866 227364 632898
rect 229686 633454 229926 633486
rect 229686 633218 229688 633454
rect 229924 633218 229926 633454
rect 229686 633134 229926 633218
rect 229686 632898 229688 633134
rect 229924 632898 229926 633134
rect 229686 632866 229926 632898
rect 230338 633454 230578 633486
rect 230338 633218 230340 633454
rect 230576 633218 230578 633454
rect 230338 633134 230578 633218
rect 230338 632898 230340 633134
rect 230576 632898 230578 633134
rect 230338 632866 230578 632898
rect 231144 633454 231384 633486
rect 231144 633218 231146 633454
rect 231382 633218 231384 633454
rect 231144 633134 231384 633218
rect 231144 632898 231146 633134
rect 231382 632898 231384 633134
rect 231144 632866 231384 632898
rect 240144 633454 240384 633486
rect 240144 633218 240146 633454
rect 240382 633218 240384 633454
rect 240144 633134 240384 633218
rect 240144 632898 240146 633134
rect 240382 632898 240384 633134
rect 240144 632866 240384 632898
rect 249144 633454 249384 633486
rect 249144 633218 249146 633454
rect 249382 633218 249384 633454
rect 249144 633134 249384 633218
rect 249144 632898 249146 633134
rect 249382 632898 249384 633134
rect 249144 632866 249384 632898
rect 258144 633454 258384 633486
rect 258144 633218 258146 633454
rect 258382 633218 258384 633454
rect 258144 633134 258384 633218
rect 258144 632898 258146 633134
rect 258382 632898 258384 633134
rect 258144 632866 258384 632898
rect 267144 633454 267384 633486
rect 267144 633218 267146 633454
rect 267382 633218 267384 633454
rect 267144 633134 267384 633218
rect 267144 632898 267146 633134
rect 267382 632898 267384 633134
rect 267144 632866 267384 632898
rect 269706 633454 269946 633486
rect 269706 633218 269708 633454
rect 269944 633218 269946 633454
rect 269706 633134 269946 633218
rect 269706 632898 269708 633134
rect 269944 632898 269946 633134
rect 269706 632866 269946 632898
rect 270358 633454 270598 633486
rect 270358 633218 270360 633454
rect 270596 633218 270598 633454
rect 270358 633134 270598 633218
rect 270358 632898 270360 633134
rect 270596 632898 270598 633134
rect 270358 632866 270598 632898
rect 271164 633454 271404 633486
rect 271164 633218 271166 633454
rect 271402 633218 271404 633454
rect 271164 633134 271404 633218
rect 271164 632898 271166 633134
rect 271402 632898 271404 633134
rect 271164 632866 271404 632898
rect 280164 633454 280404 633486
rect 280164 633218 280166 633454
rect 280402 633218 280404 633454
rect 280164 633134 280404 633218
rect 280164 632898 280166 633134
rect 280402 632898 280404 633134
rect 280164 632866 280404 632898
rect 289164 633454 289404 633486
rect 289164 633218 289166 633454
rect 289402 633218 289404 633454
rect 289164 633134 289404 633218
rect 289164 632898 289166 633134
rect 289402 632898 289404 633134
rect 289164 632866 289404 632898
rect 298164 633454 298404 633486
rect 298164 633218 298166 633454
rect 298402 633218 298404 633454
rect 298164 633134 298404 633218
rect 298164 632898 298166 633134
rect 298402 632898 298404 633134
rect 298164 632866 298404 632898
rect 307164 633454 307404 633486
rect 307164 633218 307166 633454
rect 307402 633218 307404 633454
rect 307164 633134 307404 633218
rect 307164 632898 307166 633134
rect 307402 632898 307404 633134
rect 307164 632866 307404 632898
rect 309726 633454 309966 633486
rect 309726 633218 309728 633454
rect 309964 633218 309966 633454
rect 309726 633134 309966 633218
rect 309726 632898 309728 633134
rect 309964 632898 309966 633134
rect 309726 632866 309966 632898
rect 311378 633454 311618 633486
rect 311378 633218 311380 633454
rect 311616 633218 311618 633454
rect 311378 633134 311618 633218
rect 311378 632898 311380 633134
rect 311616 632898 311618 633134
rect 311378 632866 311618 632898
rect 312184 633454 312424 633486
rect 312184 633218 312186 633454
rect 312422 633218 312424 633454
rect 312184 633134 312424 633218
rect 312184 632898 312186 633134
rect 312422 632898 312424 633134
rect 312184 632866 312424 632898
rect 321184 633454 321424 633486
rect 321184 633218 321186 633454
rect 321422 633218 321424 633454
rect 321184 633134 321424 633218
rect 321184 632898 321186 633134
rect 321422 632898 321424 633134
rect 321184 632866 321424 632898
rect 330184 633454 330424 633486
rect 330184 633218 330186 633454
rect 330422 633218 330424 633454
rect 330184 633134 330424 633218
rect 330184 632898 330186 633134
rect 330422 632898 330424 633134
rect 330184 632866 330424 632898
rect 339184 633454 339424 633486
rect 339184 633218 339186 633454
rect 339422 633218 339424 633454
rect 339184 633134 339424 633218
rect 339184 632898 339186 633134
rect 339422 632898 339424 633134
rect 339184 632866 339424 632898
rect 348184 633454 348424 633486
rect 348184 633218 348186 633454
rect 348422 633218 348424 633454
rect 348184 633134 348424 633218
rect 348184 632898 348186 633134
rect 348422 632898 348424 633134
rect 348184 632866 348424 632898
rect 350746 633454 350986 633486
rect 350746 633218 350748 633454
rect 350984 633218 350986 633454
rect 350746 633134 350986 633218
rect 350746 632898 350748 633134
rect 350984 632898 350986 633134
rect 350746 632866 350986 632898
rect 352398 633454 352638 633486
rect 352398 633218 352400 633454
rect 352636 633218 352638 633454
rect 352398 633134 352638 633218
rect 352398 632898 352400 633134
rect 352636 632898 352638 633134
rect 352398 632866 352638 632898
rect 353204 633454 353444 633486
rect 353204 633218 353206 633454
rect 353442 633218 353444 633454
rect 353204 633134 353444 633218
rect 353204 632898 353206 633134
rect 353442 632898 353444 633134
rect 353204 632866 353444 632898
rect 362204 633454 362444 633486
rect 362204 633218 362206 633454
rect 362442 633218 362444 633454
rect 362204 633134 362444 633218
rect 362204 632898 362206 633134
rect 362442 632898 362444 633134
rect 362204 632866 362444 632898
rect 371204 633454 371444 633486
rect 371204 633218 371206 633454
rect 371442 633218 371444 633454
rect 371204 633134 371444 633218
rect 371204 632898 371206 633134
rect 371442 632898 371444 633134
rect 371204 632866 371444 632898
rect 380204 633454 380444 633486
rect 380204 633218 380206 633454
rect 380442 633218 380444 633454
rect 380204 633134 380444 633218
rect 380204 632898 380206 633134
rect 380442 632898 380444 633134
rect 380204 632866 380444 632898
rect 389204 633454 389444 633486
rect 389204 633218 389206 633454
rect 389442 633218 389444 633454
rect 389204 633134 389444 633218
rect 389204 632898 389206 633134
rect 389442 632898 389444 633134
rect 389204 632866 389444 632898
rect 391766 633454 392006 633486
rect 391766 633218 391768 633454
rect 392004 633218 392006 633454
rect 391766 633134 392006 633218
rect 391766 632898 391768 633134
rect 392004 632898 392006 633134
rect 391766 632866 392006 632898
rect 392418 633454 392658 633486
rect 392418 633218 392420 633454
rect 392656 633218 392658 633454
rect 392418 633134 392658 633218
rect 392418 632898 392420 633134
rect 392656 632898 392658 633134
rect 392418 632866 392658 632898
rect 393224 633454 393464 633486
rect 393224 633218 393226 633454
rect 393462 633218 393464 633454
rect 393224 633134 393464 633218
rect 393224 632898 393226 633134
rect 393462 632898 393464 633134
rect 393224 632866 393464 632898
rect 402224 633454 402464 633486
rect 402224 633218 402226 633454
rect 402462 633218 402464 633454
rect 402224 633134 402464 633218
rect 402224 632898 402226 633134
rect 402462 632898 402464 633134
rect 402224 632866 402464 632898
rect 411224 633454 411464 633486
rect 411224 633218 411226 633454
rect 411462 633218 411464 633454
rect 411224 633134 411464 633218
rect 411224 632898 411226 633134
rect 411462 632898 411464 633134
rect 411224 632866 411464 632898
rect 420224 633454 420464 633486
rect 420224 633218 420226 633454
rect 420462 633218 420464 633454
rect 420224 633134 420464 633218
rect 420224 632898 420226 633134
rect 420462 632898 420464 633134
rect 420224 632866 420464 632898
rect 429224 633454 429464 633486
rect 429224 633218 429226 633454
rect 429462 633218 429464 633454
rect 429224 633134 429464 633218
rect 429224 632898 429226 633134
rect 429462 632898 429464 633134
rect 429224 632866 429464 632898
rect 431786 633454 432026 633486
rect 431786 633218 431788 633454
rect 432024 633218 432026 633454
rect 431786 633134 432026 633218
rect 431786 632898 431788 633134
rect 432024 632898 432026 633134
rect 431786 632866 432026 632898
rect 432438 633454 432678 633486
rect 432438 633218 432440 633454
rect 432676 633218 432678 633454
rect 432438 633134 432678 633218
rect 432438 632898 432440 633134
rect 432676 632898 432678 633134
rect 432438 632866 432678 632898
rect 433244 633454 433484 633486
rect 433244 633218 433246 633454
rect 433482 633218 433484 633454
rect 433244 633134 433484 633218
rect 433244 632898 433246 633134
rect 433482 632898 433484 633134
rect 433244 632866 433484 632898
rect 439790 633454 440030 633486
rect 439790 633218 439792 633454
rect 440028 633218 440030 633454
rect 439790 633134 440030 633218
rect 439790 632898 439792 633134
rect 440028 632898 440030 633134
rect 439790 632866 440030 632898
rect 457008 633454 457248 633486
rect 457008 633218 457010 633454
rect 457246 633218 457248 633454
rect 457008 633134 457248 633218
rect 457008 632898 457010 633134
rect 457246 632898 457248 633134
rect 457008 632866 457248 632898
rect 476596 633454 476944 633486
rect 476596 633218 476652 633454
rect 476888 633218 476944 633454
rect 476596 633134 476944 633218
rect 476596 632898 476652 633134
rect 476888 632898 476944 633134
rect 476596 632866 476944 632898
rect 571660 633454 572008 633486
rect 571660 633218 571716 633454
rect 571952 633218 572008 633454
rect 571660 633134 572008 633218
rect 571660 632898 571716 633134
rect 571952 632898 572008 633134
rect 571660 632866 572008 632898
rect 579288 633454 579888 633486
rect 579288 633218 579470 633454
rect 579706 633218 579888 633454
rect 579288 633134 579888 633218
rect 579288 632898 579470 633134
rect 579706 632898 579888 633134
rect 579288 632866 579888 632898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect 5200 615454 5800 615486
rect 5200 615218 5382 615454
rect 5618 615218 5800 615454
rect 5200 615134 5800 615218
rect 5200 614898 5382 615134
rect 5618 614898 5800 615134
rect 5200 614866 5800 614898
rect 12976 615454 13324 615486
rect 12976 615218 13032 615454
rect 13268 615218 13324 615454
rect 12976 615134 13324 615218
rect 12976 614898 13032 615134
rect 13268 614898 13324 615134
rect 12976 614866 13324 614898
rect 106680 615454 107028 615486
rect 106680 615218 106736 615454
rect 106972 615218 107028 615454
rect 106680 615134 107028 615218
rect 106680 614898 106736 615134
rect 106972 614898 107028 615134
rect 106680 614866 107028 614898
rect 127456 615454 127696 615486
rect 127456 615218 127458 615454
rect 127694 615218 127696 615454
rect 127456 615134 127696 615218
rect 127456 614898 127458 615134
rect 127694 614898 127696 615134
rect 127456 614866 127696 614898
rect 140654 615454 140894 615486
rect 140654 615218 140656 615454
rect 140892 615218 140894 615454
rect 140654 615134 140894 615218
rect 140654 614898 140656 615134
rect 140892 614898 140894 615134
rect 140654 614866 140894 614898
rect 141500 615454 141740 615486
rect 141500 615218 141502 615454
rect 141738 615218 141740 615454
rect 141500 615134 141740 615218
rect 141500 614898 141502 615134
rect 141738 614898 141740 615134
rect 141500 614866 141740 614898
rect 147286 615454 147526 615486
rect 147286 615218 147288 615454
rect 147524 615218 147526 615454
rect 147286 615134 147526 615218
rect 147286 614898 147288 615134
rect 147524 614898 147526 615134
rect 147286 614866 147526 614898
rect 149658 615454 149898 615486
rect 149658 615218 149660 615454
rect 149896 615218 149898 615454
rect 149658 615134 149898 615218
rect 149658 614898 149660 615134
rect 149896 614898 149898 615134
rect 149658 614866 149898 614898
rect 150504 615454 150744 615486
rect 150504 615218 150506 615454
rect 150742 615218 150744 615454
rect 150504 615134 150744 615218
rect 150504 614898 150506 615134
rect 150742 614898 150744 615134
rect 150504 614866 150744 614898
rect 159504 615454 159744 615486
rect 159504 615218 159506 615454
rect 159742 615218 159744 615454
rect 159504 615134 159744 615218
rect 159504 614898 159506 615134
rect 159742 614898 159744 615134
rect 159504 614866 159744 614898
rect 168504 615454 168744 615486
rect 168504 615218 168506 615454
rect 168742 615218 168744 615454
rect 168504 615134 168744 615218
rect 168504 614898 168506 615134
rect 168742 614898 168744 615134
rect 168504 614866 168744 614898
rect 177504 615454 177744 615486
rect 177504 615218 177506 615454
rect 177742 615218 177744 615454
rect 177504 615134 177744 615218
rect 177504 614898 177506 615134
rect 177742 614898 177744 615134
rect 177504 614866 177744 614898
rect 186504 615454 186744 615486
rect 186504 615218 186506 615454
rect 186742 615218 186744 615454
rect 186504 615134 186744 615218
rect 186504 614898 186506 615134
rect 186742 614898 186744 615134
rect 186504 614866 186744 614898
rect 188306 615454 188546 615486
rect 188306 615218 188308 615454
rect 188544 615218 188546 615454
rect 188306 615134 188546 615218
rect 188306 614898 188308 615134
rect 188544 614898 188546 615134
rect 188306 614866 188546 614898
rect 190678 615454 190918 615486
rect 190678 615218 190680 615454
rect 190916 615218 190918 615454
rect 190678 615134 190918 615218
rect 190678 614898 190680 615134
rect 190916 614898 190918 615134
rect 190678 614866 190918 614898
rect 191524 615454 191764 615486
rect 191524 615218 191526 615454
rect 191762 615218 191764 615454
rect 191524 615134 191764 615218
rect 191524 614898 191526 615134
rect 191762 614898 191764 615134
rect 191524 614866 191764 614898
rect 200524 615454 200764 615486
rect 200524 615218 200526 615454
rect 200762 615218 200764 615454
rect 200524 615134 200764 615218
rect 200524 614898 200526 615134
rect 200762 614898 200764 615134
rect 200524 614866 200764 614898
rect 209524 615454 209764 615486
rect 209524 615218 209526 615454
rect 209762 615218 209764 615454
rect 209524 615134 209764 615218
rect 209524 614898 209526 615134
rect 209762 614898 209764 615134
rect 209524 614866 209764 614898
rect 218524 615454 218764 615486
rect 218524 615218 218526 615454
rect 218762 615218 218764 615454
rect 218524 615134 218764 615218
rect 218524 614898 218526 615134
rect 218762 614898 218764 615134
rect 218524 614866 218764 614898
rect 227524 615454 227764 615486
rect 227524 615218 227526 615454
rect 227762 615218 227764 615454
rect 227524 615134 227764 615218
rect 227524 614898 227526 615134
rect 227762 614898 227764 615134
rect 227524 614866 227764 614898
rect 229326 615454 229566 615486
rect 229326 615218 229328 615454
rect 229564 615218 229566 615454
rect 229326 615134 229566 615218
rect 229326 614898 229328 615134
rect 229564 614898 229566 615134
rect 229326 614866 229566 614898
rect 230698 615454 230938 615486
rect 230698 615218 230700 615454
rect 230936 615218 230938 615454
rect 230698 615134 230938 615218
rect 230698 614898 230700 615134
rect 230936 614898 230938 615134
rect 230698 614866 230938 614898
rect 231544 615454 231784 615486
rect 231544 615218 231546 615454
rect 231782 615218 231784 615454
rect 231544 615134 231784 615218
rect 231544 614898 231546 615134
rect 231782 614898 231784 615134
rect 231544 614866 231784 614898
rect 240544 615454 240784 615486
rect 240544 615218 240546 615454
rect 240782 615218 240784 615454
rect 240544 615134 240784 615218
rect 240544 614898 240546 615134
rect 240782 614898 240784 615134
rect 240544 614866 240784 614898
rect 249544 615454 249784 615486
rect 249544 615218 249546 615454
rect 249782 615218 249784 615454
rect 249544 615134 249784 615218
rect 249544 614898 249546 615134
rect 249782 614898 249784 615134
rect 249544 614866 249784 614898
rect 258544 615454 258784 615486
rect 258544 615218 258546 615454
rect 258782 615218 258784 615454
rect 258544 615134 258784 615218
rect 258544 614898 258546 615134
rect 258782 614898 258784 615134
rect 258544 614866 258784 614898
rect 267544 615454 267784 615486
rect 267544 615218 267546 615454
rect 267782 615218 267784 615454
rect 267544 615134 267784 615218
rect 267544 614898 267546 615134
rect 267782 614898 267784 615134
rect 267544 614866 267784 614898
rect 269346 615454 269586 615486
rect 269346 615218 269348 615454
rect 269584 615218 269586 615454
rect 269346 615134 269586 615218
rect 269346 614898 269348 615134
rect 269584 614898 269586 615134
rect 269346 614866 269586 614898
rect 270718 615454 270958 615486
rect 270718 615218 270720 615454
rect 270956 615218 270958 615454
rect 270718 615134 270958 615218
rect 270718 614898 270720 615134
rect 270956 614898 270958 615134
rect 270718 614866 270958 614898
rect 271564 615454 271804 615486
rect 271564 615218 271566 615454
rect 271802 615218 271804 615454
rect 271564 615134 271804 615218
rect 271564 614898 271566 615134
rect 271802 614898 271804 615134
rect 271564 614866 271804 614898
rect 280564 615454 280804 615486
rect 280564 615218 280566 615454
rect 280802 615218 280804 615454
rect 280564 615134 280804 615218
rect 280564 614898 280566 615134
rect 280802 614898 280804 615134
rect 280564 614866 280804 614898
rect 289564 615454 289804 615486
rect 289564 615218 289566 615454
rect 289802 615218 289804 615454
rect 289564 615134 289804 615218
rect 289564 614898 289566 615134
rect 289802 614898 289804 615134
rect 289564 614866 289804 614898
rect 298564 615454 298804 615486
rect 298564 615218 298566 615454
rect 298802 615218 298804 615454
rect 298564 615134 298804 615218
rect 298564 614898 298566 615134
rect 298802 614898 298804 615134
rect 298564 614866 298804 614898
rect 307564 615454 307804 615486
rect 307564 615218 307566 615454
rect 307802 615218 307804 615454
rect 307564 615134 307804 615218
rect 307564 614898 307566 615134
rect 307802 614898 307804 615134
rect 307564 614866 307804 614898
rect 309366 615454 309606 615486
rect 309366 615218 309368 615454
rect 309604 615218 309606 615454
rect 309366 615134 309606 615218
rect 309366 614898 309368 615134
rect 309604 614898 309606 615134
rect 309366 614866 309606 614898
rect 311738 615454 311978 615486
rect 311738 615218 311740 615454
rect 311976 615218 311978 615454
rect 311738 615134 311978 615218
rect 311738 614898 311740 615134
rect 311976 614898 311978 615134
rect 311738 614866 311978 614898
rect 312584 615454 312824 615486
rect 312584 615218 312586 615454
rect 312822 615218 312824 615454
rect 312584 615134 312824 615218
rect 312584 614898 312586 615134
rect 312822 614898 312824 615134
rect 312584 614866 312824 614898
rect 321584 615454 321824 615486
rect 321584 615218 321586 615454
rect 321822 615218 321824 615454
rect 321584 615134 321824 615218
rect 321584 614898 321586 615134
rect 321822 614898 321824 615134
rect 321584 614866 321824 614898
rect 330584 615454 330824 615486
rect 330584 615218 330586 615454
rect 330822 615218 330824 615454
rect 330584 615134 330824 615218
rect 330584 614898 330586 615134
rect 330822 614898 330824 615134
rect 330584 614866 330824 614898
rect 339584 615454 339824 615486
rect 339584 615218 339586 615454
rect 339822 615218 339824 615454
rect 339584 615134 339824 615218
rect 339584 614898 339586 615134
rect 339822 614898 339824 615134
rect 339584 614866 339824 614898
rect 348584 615454 348824 615486
rect 348584 615218 348586 615454
rect 348822 615218 348824 615454
rect 348584 615134 348824 615218
rect 348584 614898 348586 615134
rect 348822 614898 348824 615134
rect 348584 614866 348824 614898
rect 350386 615454 350626 615486
rect 350386 615218 350388 615454
rect 350624 615218 350626 615454
rect 350386 615134 350626 615218
rect 350386 614898 350388 615134
rect 350624 614898 350626 615134
rect 350386 614866 350626 614898
rect 352758 615454 352998 615486
rect 352758 615218 352760 615454
rect 352996 615218 352998 615454
rect 352758 615134 352998 615218
rect 352758 614898 352760 615134
rect 352996 614898 352998 615134
rect 352758 614866 352998 614898
rect 353604 615454 353844 615486
rect 353604 615218 353606 615454
rect 353842 615218 353844 615454
rect 353604 615134 353844 615218
rect 353604 614898 353606 615134
rect 353842 614898 353844 615134
rect 353604 614866 353844 614898
rect 362604 615454 362844 615486
rect 362604 615218 362606 615454
rect 362842 615218 362844 615454
rect 362604 615134 362844 615218
rect 362604 614898 362606 615134
rect 362842 614898 362844 615134
rect 362604 614866 362844 614898
rect 371604 615454 371844 615486
rect 371604 615218 371606 615454
rect 371842 615218 371844 615454
rect 371604 615134 371844 615218
rect 371604 614898 371606 615134
rect 371842 614898 371844 615134
rect 371604 614866 371844 614898
rect 380604 615454 380844 615486
rect 380604 615218 380606 615454
rect 380842 615218 380844 615454
rect 380604 615134 380844 615218
rect 380604 614898 380606 615134
rect 380842 614898 380844 615134
rect 380604 614866 380844 614898
rect 389604 615454 389844 615486
rect 389604 615218 389606 615454
rect 389842 615218 389844 615454
rect 389604 615134 389844 615218
rect 389604 614898 389606 615134
rect 389842 614898 389844 615134
rect 389604 614866 389844 614898
rect 391406 615454 391646 615486
rect 391406 615218 391408 615454
rect 391644 615218 391646 615454
rect 391406 615134 391646 615218
rect 391406 614898 391408 615134
rect 391644 614898 391646 615134
rect 391406 614866 391646 614898
rect 392778 615454 393018 615486
rect 392778 615218 392780 615454
rect 393016 615218 393018 615454
rect 392778 615134 393018 615218
rect 392778 614898 392780 615134
rect 393016 614898 393018 615134
rect 392778 614866 393018 614898
rect 393624 615454 393864 615486
rect 393624 615218 393626 615454
rect 393862 615218 393864 615454
rect 393624 615134 393864 615218
rect 393624 614898 393626 615134
rect 393862 614898 393864 615134
rect 393624 614866 393864 614898
rect 402624 615454 402864 615486
rect 402624 615218 402626 615454
rect 402862 615218 402864 615454
rect 402624 615134 402864 615218
rect 402624 614898 402626 615134
rect 402862 614898 402864 615134
rect 402624 614866 402864 614898
rect 411624 615454 411864 615486
rect 411624 615218 411626 615454
rect 411862 615218 411864 615454
rect 411624 615134 411864 615218
rect 411624 614898 411626 615134
rect 411862 614898 411864 615134
rect 411624 614866 411864 614898
rect 420624 615454 420864 615486
rect 420624 615218 420626 615454
rect 420862 615218 420864 615454
rect 420624 615134 420864 615218
rect 420624 614898 420626 615134
rect 420862 614898 420864 615134
rect 420624 614866 420864 614898
rect 429624 615454 429864 615486
rect 429624 615218 429626 615454
rect 429862 615218 429864 615454
rect 429624 615134 429864 615218
rect 429624 614898 429626 615134
rect 429862 614898 429864 615134
rect 429624 614866 429864 614898
rect 431426 615454 431666 615486
rect 431426 615218 431428 615454
rect 431664 615218 431666 615454
rect 431426 615134 431666 615218
rect 431426 614898 431428 615134
rect 431664 614898 431666 615134
rect 431426 614866 431666 614898
rect 432798 615454 433038 615486
rect 432798 615218 432800 615454
rect 433036 615218 433038 615454
rect 432798 615134 433038 615218
rect 432798 614898 432800 615134
rect 433036 614898 433038 615134
rect 432798 614866 433038 614898
rect 433644 615454 433884 615486
rect 433644 615218 433646 615454
rect 433882 615218 433884 615454
rect 433644 615134 433884 615218
rect 433644 614898 433646 615134
rect 433882 614898 433884 615134
rect 433644 614866 433884 614898
rect 439430 615454 439670 615486
rect 439430 615218 439432 615454
rect 439668 615218 439670 615454
rect 439430 615134 439670 615218
rect 439430 614898 439432 615134
rect 439668 614898 439670 615134
rect 439430 614866 439670 614898
rect 456608 615454 456848 615486
rect 456608 615218 456610 615454
rect 456846 615218 456848 615454
rect 456608 615134 456848 615218
rect 456608 614898 456610 615134
rect 456846 614898 456848 615134
rect 456608 614866 456848 614898
rect 477276 615454 477624 615486
rect 477276 615218 477332 615454
rect 477568 615218 477624 615454
rect 477276 615134 477624 615218
rect 477276 614898 477332 615134
rect 477568 614898 477624 615134
rect 477276 614866 477624 614898
rect 570980 615454 571328 615486
rect 570980 615218 571036 615454
rect 571272 615218 571328 615454
rect 570980 615134 571328 615218
rect 570980 614898 571036 615134
rect 571272 614898 571328 615134
rect 570980 614866 571328 614898
rect 578488 615454 579088 615486
rect 578488 615218 578670 615454
rect 578906 615218 579088 615454
rect 578488 615134 579088 615218
rect 578488 614898 578670 615134
rect 578906 614898 579088 615134
rect 578488 614866 579088 614898
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 4400 597454 5000 597486
rect 4400 597218 4582 597454
rect 4818 597218 5000 597454
rect 4400 597134 5000 597218
rect 4400 596898 4582 597134
rect 4818 596898 5000 597134
rect 4400 596866 5000 596898
rect 12296 597454 12644 597486
rect 12296 597218 12352 597454
rect 12588 597218 12644 597454
rect 12296 597134 12644 597218
rect 12296 596898 12352 597134
rect 12588 596898 12644 597134
rect 12296 596866 12644 596898
rect 107360 597454 107708 597486
rect 107360 597218 107416 597454
rect 107652 597218 107708 597454
rect 107360 597134 107708 597218
rect 107360 596898 107416 597134
rect 107652 596898 107708 597134
rect 107360 596866 107708 596898
rect 127056 597454 127296 597486
rect 127056 597218 127058 597454
rect 127294 597218 127296 597454
rect 127056 597134 127296 597218
rect 127056 596898 127058 597134
rect 127294 596898 127296 597134
rect 127056 596866 127296 596898
rect 140294 597454 140534 597486
rect 140294 597218 140296 597454
rect 140532 597218 140534 597454
rect 140294 597134 140534 597218
rect 140294 596898 140296 597134
rect 140532 596898 140534 597134
rect 140294 596866 140534 596898
rect 141100 597454 141340 597486
rect 141100 597218 141102 597454
rect 141338 597218 141340 597454
rect 141100 597134 141340 597218
rect 141100 596898 141102 597134
rect 141338 596898 141340 597134
rect 141100 596866 141340 596898
rect 147646 597454 147886 597486
rect 147646 597218 147648 597454
rect 147884 597218 147886 597454
rect 147646 597134 147886 597218
rect 147646 596898 147648 597134
rect 147884 596898 147886 597134
rect 147646 596866 147886 596898
rect 149298 597454 149538 597486
rect 149298 597218 149300 597454
rect 149536 597218 149538 597454
rect 149298 597134 149538 597218
rect 149298 596898 149300 597134
rect 149536 596898 149538 597134
rect 149298 596866 149538 596898
rect 150104 597454 150344 597486
rect 150104 597218 150106 597454
rect 150342 597218 150344 597454
rect 150104 597134 150344 597218
rect 150104 596898 150106 597134
rect 150342 596898 150344 597134
rect 150104 596866 150344 596898
rect 159104 597454 159344 597486
rect 159104 597218 159106 597454
rect 159342 597218 159344 597454
rect 159104 597134 159344 597218
rect 159104 596898 159106 597134
rect 159342 596898 159344 597134
rect 159104 596866 159344 596898
rect 168104 597454 168344 597486
rect 168104 597218 168106 597454
rect 168342 597218 168344 597454
rect 168104 597134 168344 597218
rect 168104 596898 168106 597134
rect 168342 596898 168344 597134
rect 168104 596866 168344 596898
rect 177104 597454 177344 597486
rect 177104 597218 177106 597454
rect 177342 597218 177344 597454
rect 177104 597134 177344 597218
rect 177104 596898 177106 597134
rect 177342 596898 177344 597134
rect 177104 596866 177344 596898
rect 186104 597454 186344 597486
rect 186104 597218 186106 597454
rect 186342 597218 186344 597454
rect 186104 597134 186344 597218
rect 186104 596898 186106 597134
rect 186342 596898 186344 597134
rect 186104 596866 186344 596898
rect 188666 597454 188906 597486
rect 188666 597218 188668 597454
rect 188904 597218 188906 597454
rect 188666 597134 188906 597218
rect 188666 596898 188668 597134
rect 188904 596898 188906 597134
rect 188666 596866 188906 596898
rect 189766 597454 190006 597486
rect 189766 597218 189768 597454
rect 190004 597218 190006 597454
rect 189766 597134 190006 597218
rect 189766 596898 189768 597134
rect 190004 596898 190006 597134
rect 189766 596866 190006 596898
rect 190318 597454 190558 597486
rect 190318 597218 190320 597454
rect 190556 597218 190558 597454
rect 190318 597134 190558 597218
rect 190318 596898 190320 597134
rect 190556 596898 190558 597134
rect 190318 596866 190558 596898
rect 191124 597454 191364 597486
rect 191124 597218 191126 597454
rect 191362 597218 191364 597454
rect 191124 597134 191364 597218
rect 191124 596898 191126 597134
rect 191362 596898 191364 597134
rect 191124 596866 191364 596898
rect 200124 597454 200364 597486
rect 200124 597218 200126 597454
rect 200362 597218 200364 597454
rect 200124 597134 200364 597218
rect 200124 596898 200126 597134
rect 200362 596898 200364 597134
rect 200124 596866 200364 596898
rect 209124 597454 209364 597486
rect 209124 597218 209126 597454
rect 209362 597218 209364 597454
rect 209124 597134 209364 597218
rect 209124 596898 209126 597134
rect 209362 596898 209364 597134
rect 209124 596866 209364 596898
rect 218124 597454 218364 597486
rect 218124 597218 218126 597454
rect 218362 597218 218364 597454
rect 218124 597134 218364 597218
rect 218124 596898 218126 597134
rect 218362 596898 218364 597134
rect 218124 596866 218364 596898
rect 227124 597454 227364 597486
rect 227124 597218 227126 597454
rect 227362 597218 227364 597454
rect 227124 597134 227364 597218
rect 227124 596898 227126 597134
rect 227362 596898 227364 597134
rect 227124 596866 227364 596898
rect 229686 597454 229926 597486
rect 229686 597218 229688 597454
rect 229924 597218 229926 597454
rect 229686 597134 229926 597218
rect 229686 596898 229688 597134
rect 229924 596898 229926 597134
rect 229686 596866 229926 596898
rect 230338 597454 230578 597486
rect 230338 597218 230340 597454
rect 230576 597218 230578 597454
rect 230338 597134 230578 597218
rect 230338 596898 230340 597134
rect 230576 596898 230578 597134
rect 230338 596866 230578 596898
rect 231144 597454 231384 597486
rect 231144 597218 231146 597454
rect 231382 597218 231384 597454
rect 231144 597134 231384 597218
rect 231144 596898 231146 597134
rect 231382 596898 231384 597134
rect 231144 596866 231384 596898
rect 240144 597454 240384 597486
rect 240144 597218 240146 597454
rect 240382 597218 240384 597454
rect 240144 597134 240384 597218
rect 240144 596898 240146 597134
rect 240382 596898 240384 597134
rect 240144 596866 240384 596898
rect 249144 597454 249384 597486
rect 249144 597218 249146 597454
rect 249382 597218 249384 597454
rect 249144 597134 249384 597218
rect 249144 596898 249146 597134
rect 249382 596898 249384 597134
rect 249144 596866 249384 596898
rect 258144 597454 258384 597486
rect 258144 597218 258146 597454
rect 258382 597218 258384 597454
rect 258144 597134 258384 597218
rect 258144 596898 258146 597134
rect 258382 596898 258384 597134
rect 258144 596866 258384 596898
rect 267144 597454 267384 597486
rect 267144 597218 267146 597454
rect 267382 597218 267384 597454
rect 267144 597134 267384 597218
rect 267144 596898 267146 597134
rect 267382 596898 267384 597134
rect 267144 596866 267384 596898
rect 269706 597454 269946 597486
rect 269706 597218 269708 597454
rect 269944 597218 269946 597454
rect 269706 597134 269946 597218
rect 269706 596898 269708 597134
rect 269944 596898 269946 597134
rect 269706 596866 269946 596898
rect 270358 597454 270598 597486
rect 270358 597218 270360 597454
rect 270596 597218 270598 597454
rect 270358 597134 270598 597218
rect 270358 596898 270360 597134
rect 270596 596898 270598 597134
rect 270358 596866 270598 596898
rect 271164 597454 271404 597486
rect 271164 597218 271166 597454
rect 271402 597218 271404 597454
rect 271164 597134 271404 597218
rect 271164 596898 271166 597134
rect 271402 596898 271404 597134
rect 271164 596866 271404 596898
rect 280164 597454 280404 597486
rect 280164 597218 280166 597454
rect 280402 597218 280404 597454
rect 280164 597134 280404 597218
rect 280164 596898 280166 597134
rect 280402 596898 280404 597134
rect 280164 596866 280404 596898
rect 289164 597454 289404 597486
rect 289164 597218 289166 597454
rect 289402 597218 289404 597454
rect 289164 597134 289404 597218
rect 289164 596898 289166 597134
rect 289402 596898 289404 597134
rect 289164 596866 289404 596898
rect 298164 597454 298404 597486
rect 298164 597218 298166 597454
rect 298402 597218 298404 597454
rect 298164 597134 298404 597218
rect 298164 596898 298166 597134
rect 298402 596898 298404 597134
rect 298164 596866 298404 596898
rect 307164 597454 307404 597486
rect 307164 597218 307166 597454
rect 307402 597218 307404 597454
rect 307164 597134 307404 597218
rect 307164 596898 307166 597134
rect 307402 596898 307404 597134
rect 307164 596866 307404 596898
rect 309726 597454 309966 597486
rect 309726 597218 309728 597454
rect 309964 597218 309966 597454
rect 309726 597134 309966 597218
rect 309726 596898 309728 597134
rect 309964 596898 309966 597134
rect 309726 596866 309966 596898
rect 311378 597454 311618 597486
rect 311378 597218 311380 597454
rect 311616 597218 311618 597454
rect 311378 597134 311618 597218
rect 311378 596898 311380 597134
rect 311616 596898 311618 597134
rect 311378 596866 311618 596898
rect 312184 597454 312424 597486
rect 312184 597218 312186 597454
rect 312422 597218 312424 597454
rect 312184 597134 312424 597218
rect 312184 596898 312186 597134
rect 312422 596898 312424 597134
rect 312184 596866 312424 596898
rect 321184 597454 321424 597486
rect 321184 597218 321186 597454
rect 321422 597218 321424 597454
rect 321184 597134 321424 597218
rect 321184 596898 321186 597134
rect 321422 596898 321424 597134
rect 321184 596866 321424 596898
rect 330184 597454 330424 597486
rect 330184 597218 330186 597454
rect 330422 597218 330424 597454
rect 330184 597134 330424 597218
rect 330184 596898 330186 597134
rect 330422 596898 330424 597134
rect 330184 596866 330424 596898
rect 339184 597454 339424 597486
rect 339184 597218 339186 597454
rect 339422 597218 339424 597454
rect 339184 597134 339424 597218
rect 339184 596898 339186 597134
rect 339422 596898 339424 597134
rect 339184 596866 339424 596898
rect 348184 597454 348424 597486
rect 348184 597218 348186 597454
rect 348422 597218 348424 597454
rect 348184 597134 348424 597218
rect 348184 596898 348186 597134
rect 348422 596898 348424 597134
rect 348184 596866 348424 596898
rect 350746 597454 350986 597486
rect 350746 597218 350748 597454
rect 350984 597218 350986 597454
rect 350746 597134 350986 597218
rect 350746 596898 350748 597134
rect 350984 596898 350986 597134
rect 350746 596866 350986 596898
rect 352398 597454 352638 597486
rect 352398 597218 352400 597454
rect 352636 597218 352638 597454
rect 352398 597134 352638 597218
rect 352398 596898 352400 597134
rect 352636 596898 352638 597134
rect 352398 596866 352638 596898
rect 353204 597454 353444 597486
rect 353204 597218 353206 597454
rect 353442 597218 353444 597454
rect 353204 597134 353444 597218
rect 353204 596898 353206 597134
rect 353442 596898 353444 597134
rect 353204 596866 353444 596898
rect 362204 597454 362444 597486
rect 362204 597218 362206 597454
rect 362442 597218 362444 597454
rect 362204 597134 362444 597218
rect 362204 596898 362206 597134
rect 362442 596898 362444 597134
rect 362204 596866 362444 596898
rect 371204 597454 371444 597486
rect 371204 597218 371206 597454
rect 371442 597218 371444 597454
rect 371204 597134 371444 597218
rect 371204 596898 371206 597134
rect 371442 596898 371444 597134
rect 371204 596866 371444 596898
rect 380204 597454 380444 597486
rect 380204 597218 380206 597454
rect 380442 597218 380444 597454
rect 380204 597134 380444 597218
rect 380204 596898 380206 597134
rect 380442 596898 380444 597134
rect 380204 596866 380444 596898
rect 389204 597454 389444 597486
rect 389204 597218 389206 597454
rect 389442 597218 389444 597454
rect 389204 597134 389444 597218
rect 389204 596898 389206 597134
rect 389442 596898 389444 597134
rect 389204 596866 389444 596898
rect 391766 597454 392006 597486
rect 391766 597218 391768 597454
rect 392004 597218 392006 597454
rect 391766 597134 392006 597218
rect 391766 596898 391768 597134
rect 392004 596898 392006 597134
rect 391766 596866 392006 596898
rect 392418 597454 392658 597486
rect 392418 597218 392420 597454
rect 392656 597218 392658 597454
rect 392418 597134 392658 597218
rect 392418 596898 392420 597134
rect 392656 596898 392658 597134
rect 392418 596866 392658 596898
rect 393224 597454 393464 597486
rect 393224 597218 393226 597454
rect 393462 597218 393464 597454
rect 393224 597134 393464 597218
rect 393224 596898 393226 597134
rect 393462 596898 393464 597134
rect 393224 596866 393464 596898
rect 402224 597454 402464 597486
rect 402224 597218 402226 597454
rect 402462 597218 402464 597454
rect 402224 597134 402464 597218
rect 402224 596898 402226 597134
rect 402462 596898 402464 597134
rect 402224 596866 402464 596898
rect 411224 597454 411464 597486
rect 411224 597218 411226 597454
rect 411462 597218 411464 597454
rect 411224 597134 411464 597218
rect 411224 596898 411226 597134
rect 411462 596898 411464 597134
rect 411224 596866 411464 596898
rect 420224 597454 420464 597486
rect 420224 597218 420226 597454
rect 420462 597218 420464 597454
rect 420224 597134 420464 597218
rect 420224 596898 420226 597134
rect 420462 596898 420464 597134
rect 420224 596866 420464 596898
rect 429224 597454 429464 597486
rect 429224 597218 429226 597454
rect 429462 597218 429464 597454
rect 429224 597134 429464 597218
rect 429224 596898 429226 597134
rect 429462 596898 429464 597134
rect 429224 596866 429464 596898
rect 431786 597454 432026 597486
rect 431786 597218 431788 597454
rect 432024 597218 432026 597454
rect 431786 597134 432026 597218
rect 431786 596898 431788 597134
rect 432024 596898 432026 597134
rect 431786 596866 432026 596898
rect 432438 597454 432678 597486
rect 432438 597218 432440 597454
rect 432676 597218 432678 597454
rect 432438 597134 432678 597218
rect 432438 596898 432440 597134
rect 432676 596898 432678 597134
rect 432438 596866 432678 596898
rect 433244 597454 433484 597486
rect 433244 597218 433246 597454
rect 433482 597218 433484 597454
rect 433244 597134 433484 597218
rect 433244 596898 433246 597134
rect 433482 596898 433484 597134
rect 433244 596866 433484 596898
rect 439790 597454 440030 597486
rect 439790 597218 439792 597454
rect 440028 597218 440030 597454
rect 439790 597134 440030 597218
rect 439790 596898 439792 597134
rect 440028 596898 440030 597134
rect 439790 596866 440030 596898
rect 457008 597454 457248 597486
rect 457008 597218 457010 597454
rect 457246 597218 457248 597454
rect 457008 597134 457248 597218
rect 457008 596898 457010 597134
rect 457246 596898 457248 597134
rect 457008 596866 457248 596898
rect 476596 597454 476944 597486
rect 476596 597218 476652 597454
rect 476888 597218 476944 597454
rect 476596 597134 476944 597218
rect 476596 596898 476652 597134
rect 476888 596898 476944 597134
rect 476596 596866 476944 596898
rect 571660 597454 572008 597486
rect 571660 597218 571716 597454
rect 571952 597218 572008 597454
rect 571660 597134 572008 597218
rect 571660 596898 571716 597134
rect 571952 596898 572008 597134
rect 571660 596866 572008 596898
rect 579288 597454 579888 597486
rect 579288 597218 579470 597454
rect 579706 597218 579888 597454
rect 579288 597134 579888 597218
rect 579288 596898 579470 597134
rect 579706 596898 579888 597134
rect 579288 596866 579888 596898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect 5200 579454 5800 579486
rect 5200 579218 5382 579454
rect 5618 579218 5800 579454
rect 5200 579134 5800 579218
rect 5200 578898 5382 579134
rect 5618 578898 5800 579134
rect 5200 578866 5800 578898
rect 12976 579454 13324 579486
rect 12976 579218 13032 579454
rect 13268 579218 13324 579454
rect 12976 579134 13324 579218
rect 12976 578898 13032 579134
rect 13268 578898 13324 579134
rect 12976 578866 13324 578898
rect 106680 579454 107028 579486
rect 106680 579218 106736 579454
rect 106972 579218 107028 579454
rect 106680 579134 107028 579218
rect 106680 578898 106736 579134
rect 106972 578898 107028 579134
rect 106680 578866 107028 578898
rect 127456 579454 127696 579486
rect 127456 579218 127458 579454
rect 127694 579218 127696 579454
rect 127456 579134 127696 579218
rect 127456 578898 127458 579134
rect 127694 578898 127696 579134
rect 127456 578866 127696 578898
rect 140654 579454 140894 579486
rect 140654 579218 140656 579454
rect 140892 579218 140894 579454
rect 140654 579134 140894 579218
rect 140654 578898 140656 579134
rect 140892 578898 140894 579134
rect 140654 578866 140894 578898
rect 141500 579454 141740 579486
rect 141500 579218 141502 579454
rect 141738 579218 141740 579454
rect 141500 579134 141740 579218
rect 141500 578898 141502 579134
rect 141738 578898 141740 579134
rect 141500 578866 141740 578898
rect 147286 579454 147526 579486
rect 147286 579218 147288 579454
rect 147524 579218 147526 579454
rect 147286 579134 147526 579218
rect 147286 578898 147288 579134
rect 147524 578898 147526 579134
rect 147286 578866 147526 578898
rect 149658 579454 149898 579486
rect 149658 579218 149660 579454
rect 149896 579218 149898 579454
rect 149658 579134 149898 579218
rect 149658 578898 149660 579134
rect 149896 578898 149898 579134
rect 149658 578866 149898 578898
rect 150504 579454 150744 579486
rect 150504 579218 150506 579454
rect 150742 579218 150744 579454
rect 150504 579134 150744 579218
rect 150504 578898 150506 579134
rect 150742 578898 150744 579134
rect 150504 578866 150744 578898
rect 159504 579454 159744 579486
rect 159504 579218 159506 579454
rect 159742 579218 159744 579454
rect 159504 579134 159744 579218
rect 159504 578898 159506 579134
rect 159742 578898 159744 579134
rect 159504 578866 159744 578898
rect 168504 579454 168744 579486
rect 168504 579218 168506 579454
rect 168742 579218 168744 579454
rect 168504 579134 168744 579218
rect 168504 578898 168506 579134
rect 168742 578898 168744 579134
rect 168504 578866 168744 578898
rect 177504 579454 177744 579486
rect 177504 579218 177506 579454
rect 177742 579218 177744 579454
rect 177504 579134 177744 579218
rect 177504 578898 177506 579134
rect 177742 578898 177744 579134
rect 177504 578866 177744 578898
rect 186504 579454 186744 579486
rect 186504 579218 186506 579454
rect 186742 579218 186744 579454
rect 186504 579134 186744 579218
rect 186504 578898 186506 579134
rect 186742 578898 186744 579134
rect 186504 578866 186744 578898
rect 188306 579454 188546 579486
rect 188306 579218 188308 579454
rect 188544 579218 188546 579454
rect 188306 579134 188546 579218
rect 188306 578898 188308 579134
rect 188544 578898 188546 579134
rect 188306 578866 188546 578898
rect 190678 579454 190918 579486
rect 190678 579218 190680 579454
rect 190916 579218 190918 579454
rect 190678 579134 190918 579218
rect 190678 578898 190680 579134
rect 190916 578898 190918 579134
rect 190678 578866 190918 578898
rect 191524 579454 191764 579486
rect 191524 579218 191526 579454
rect 191762 579218 191764 579454
rect 191524 579134 191764 579218
rect 191524 578898 191526 579134
rect 191762 578898 191764 579134
rect 191524 578866 191764 578898
rect 200524 579454 200764 579486
rect 200524 579218 200526 579454
rect 200762 579218 200764 579454
rect 200524 579134 200764 579218
rect 200524 578898 200526 579134
rect 200762 578898 200764 579134
rect 200524 578866 200764 578898
rect 209524 579454 209764 579486
rect 209524 579218 209526 579454
rect 209762 579218 209764 579454
rect 209524 579134 209764 579218
rect 209524 578898 209526 579134
rect 209762 578898 209764 579134
rect 209524 578866 209764 578898
rect 218524 579454 218764 579486
rect 218524 579218 218526 579454
rect 218762 579218 218764 579454
rect 218524 579134 218764 579218
rect 218524 578898 218526 579134
rect 218762 578898 218764 579134
rect 218524 578866 218764 578898
rect 227524 579454 227764 579486
rect 227524 579218 227526 579454
rect 227762 579218 227764 579454
rect 227524 579134 227764 579218
rect 227524 578898 227526 579134
rect 227762 578898 227764 579134
rect 227524 578866 227764 578898
rect 229326 579454 229566 579486
rect 229326 579218 229328 579454
rect 229564 579218 229566 579454
rect 229326 579134 229566 579218
rect 229326 578898 229328 579134
rect 229564 578898 229566 579134
rect 229326 578866 229566 578898
rect 230698 579454 230938 579486
rect 230698 579218 230700 579454
rect 230936 579218 230938 579454
rect 230698 579134 230938 579218
rect 230698 578898 230700 579134
rect 230936 578898 230938 579134
rect 230698 578866 230938 578898
rect 231544 579454 231784 579486
rect 231544 579218 231546 579454
rect 231782 579218 231784 579454
rect 231544 579134 231784 579218
rect 231544 578898 231546 579134
rect 231782 578898 231784 579134
rect 231544 578866 231784 578898
rect 240544 579454 240784 579486
rect 240544 579218 240546 579454
rect 240782 579218 240784 579454
rect 240544 579134 240784 579218
rect 240544 578898 240546 579134
rect 240782 578898 240784 579134
rect 240544 578866 240784 578898
rect 249544 579454 249784 579486
rect 249544 579218 249546 579454
rect 249782 579218 249784 579454
rect 249544 579134 249784 579218
rect 249544 578898 249546 579134
rect 249782 578898 249784 579134
rect 249544 578866 249784 578898
rect 258544 579454 258784 579486
rect 258544 579218 258546 579454
rect 258782 579218 258784 579454
rect 258544 579134 258784 579218
rect 258544 578898 258546 579134
rect 258782 578898 258784 579134
rect 258544 578866 258784 578898
rect 267544 579454 267784 579486
rect 267544 579218 267546 579454
rect 267782 579218 267784 579454
rect 267544 579134 267784 579218
rect 267544 578898 267546 579134
rect 267782 578898 267784 579134
rect 267544 578866 267784 578898
rect 269346 579454 269586 579486
rect 269346 579218 269348 579454
rect 269584 579218 269586 579454
rect 269346 579134 269586 579218
rect 269346 578898 269348 579134
rect 269584 578898 269586 579134
rect 269346 578866 269586 578898
rect 270718 579454 270958 579486
rect 270718 579218 270720 579454
rect 270956 579218 270958 579454
rect 270718 579134 270958 579218
rect 270718 578898 270720 579134
rect 270956 578898 270958 579134
rect 270718 578866 270958 578898
rect 271564 579454 271804 579486
rect 271564 579218 271566 579454
rect 271802 579218 271804 579454
rect 271564 579134 271804 579218
rect 271564 578898 271566 579134
rect 271802 578898 271804 579134
rect 271564 578866 271804 578898
rect 280564 579454 280804 579486
rect 280564 579218 280566 579454
rect 280802 579218 280804 579454
rect 280564 579134 280804 579218
rect 280564 578898 280566 579134
rect 280802 578898 280804 579134
rect 280564 578866 280804 578898
rect 289564 579454 289804 579486
rect 289564 579218 289566 579454
rect 289802 579218 289804 579454
rect 289564 579134 289804 579218
rect 289564 578898 289566 579134
rect 289802 578898 289804 579134
rect 289564 578866 289804 578898
rect 298564 579454 298804 579486
rect 298564 579218 298566 579454
rect 298802 579218 298804 579454
rect 298564 579134 298804 579218
rect 298564 578898 298566 579134
rect 298802 578898 298804 579134
rect 298564 578866 298804 578898
rect 307564 579454 307804 579486
rect 307564 579218 307566 579454
rect 307802 579218 307804 579454
rect 307564 579134 307804 579218
rect 307564 578898 307566 579134
rect 307802 578898 307804 579134
rect 307564 578866 307804 578898
rect 309366 579454 309606 579486
rect 309366 579218 309368 579454
rect 309604 579218 309606 579454
rect 309366 579134 309606 579218
rect 309366 578898 309368 579134
rect 309604 578898 309606 579134
rect 309366 578866 309606 578898
rect 311738 579454 311978 579486
rect 311738 579218 311740 579454
rect 311976 579218 311978 579454
rect 311738 579134 311978 579218
rect 311738 578898 311740 579134
rect 311976 578898 311978 579134
rect 311738 578866 311978 578898
rect 312584 579454 312824 579486
rect 312584 579218 312586 579454
rect 312822 579218 312824 579454
rect 312584 579134 312824 579218
rect 312584 578898 312586 579134
rect 312822 578898 312824 579134
rect 312584 578866 312824 578898
rect 321584 579454 321824 579486
rect 321584 579218 321586 579454
rect 321822 579218 321824 579454
rect 321584 579134 321824 579218
rect 321584 578898 321586 579134
rect 321822 578898 321824 579134
rect 321584 578866 321824 578898
rect 330584 579454 330824 579486
rect 330584 579218 330586 579454
rect 330822 579218 330824 579454
rect 330584 579134 330824 579218
rect 330584 578898 330586 579134
rect 330822 578898 330824 579134
rect 330584 578866 330824 578898
rect 339584 579454 339824 579486
rect 339584 579218 339586 579454
rect 339822 579218 339824 579454
rect 339584 579134 339824 579218
rect 339584 578898 339586 579134
rect 339822 578898 339824 579134
rect 339584 578866 339824 578898
rect 348584 579454 348824 579486
rect 348584 579218 348586 579454
rect 348822 579218 348824 579454
rect 348584 579134 348824 579218
rect 348584 578898 348586 579134
rect 348822 578898 348824 579134
rect 348584 578866 348824 578898
rect 350386 579454 350626 579486
rect 350386 579218 350388 579454
rect 350624 579218 350626 579454
rect 350386 579134 350626 579218
rect 350386 578898 350388 579134
rect 350624 578898 350626 579134
rect 350386 578866 350626 578898
rect 352758 579454 352998 579486
rect 352758 579218 352760 579454
rect 352996 579218 352998 579454
rect 352758 579134 352998 579218
rect 352758 578898 352760 579134
rect 352996 578898 352998 579134
rect 352758 578866 352998 578898
rect 353604 579454 353844 579486
rect 353604 579218 353606 579454
rect 353842 579218 353844 579454
rect 353604 579134 353844 579218
rect 353604 578898 353606 579134
rect 353842 578898 353844 579134
rect 353604 578866 353844 578898
rect 362604 579454 362844 579486
rect 362604 579218 362606 579454
rect 362842 579218 362844 579454
rect 362604 579134 362844 579218
rect 362604 578898 362606 579134
rect 362842 578898 362844 579134
rect 362604 578866 362844 578898
rect 371604 579454 371844 579486
rect 371604 579218 371606 579454
rect 371842 579218 371844 579454
rect 371604 579134 371844 579218
rect 371604 578898 371606 579134
rect 371842 578898 371844 579134
rect 371604 578866 371844 578898
rect 380604 579454 380844 579486
rect 380604 579218 380606 579454
rect 380842 579218 380844 579454
rect 380604 579134 380844 579218
rect 380604 578898 380606 579134
rect 380842 578898 380844 579134
rect 380604 578866 380844 578898
rect 389604 579454 389844 579486
rect 389604 579218 389606 579454
rect 389842 579218 389844 579454
rect 389604 579134 389844 579218
rect 389604 578898 389606 579134
rect 389842 578898 389844 579134
rect 389604 578866 389844 578898
rect 391406 579454 391646 579486
rect 391406 579218 391408 579454
rect 391644 579218 391646 579454
rect 391406 579134 391646 579218
rect 391406 578898 391408 579134
rect 391644 578898 391646 579134
rect 391406 578866 391646 578898
rect 392778 579454 393018 579486
rect 392778 579218 392780 579454
rect 393016 579218 393018 579454
rect 392778 579134 393018 579218
rect 392778 578898 392780 579134
rect 393016 578898 393018 579134
rect 392778 578866 393018 578898
rect 393624 579454 393864 579486
rect 393624 579218 393626 579454
rect 393862 579218 393864 579454
rect 393624 579134 393864 579218
rect 393624 578898 393626 579134
rect 393862 578898 393864 579134
rect 393624 578866 393864 578898
rect 402624 579454 402864 579486
rect 402624 579218 402626 579454
rect 402862 579218 402864 579454
rect 402624 579134 402864 579218
rect 402624 578898 402626 579134
rect 402862 578898 402864 579134
rect 402624 578866 402864 578898
rect 411624 579454 411864 579486
rect 411624 579218 411626 579454
rect 411862 579218 411864 579454
rect 411624 579134 411864 579218
rect 411624 578898 411626 579134
rect 411862 578898 411864 579134
rect 411624 578866 411864 578898
rect 420624 579454 420864 579486
rect 420624 579218 420626 579454
rect 420862 579218 420864 579454
rect 420624 579134 420864 579218
rect 420624 578898 420626 579134
rect 420862 578898 420864 579134
rect 420624 578866 420864 578898
rect 429624 579454 429864 579486
rect 429624 579218 429626 579454
rect 429862 579218 429864 579454
rect 429624 579134 429864 579218
rect 429624 578898 429626 579134
rect 429862 578898 429864 579134
rect 429624 578866 429864 578898
rect 431426 579454 431666 579486
rect 431426 579218 431428 579454
rect 431664 579218 431666 579454
rect 431426 579134 431666 579218
rect 431426 578898 431428 579134
rect 431664 578898 431666 579134
rect 431426 578866 431666 578898
rect 432798 579454 433038 579486
rect 432798 579218 432800 579454
rect 433036 579218 433038 579454
rect 432798 579134 433038 579218
rect 432798 578898 432800 579134
rect 433036 578898 433038 579134
rect 432798 578866 433038 578898
rect 433644 579454 433884 579486
rect 433644 579218 433646 579454
rect 433882 579218 433884 579454
rect 433644 579134 433884 579218
rect 433644 578898 433646 579134
rect 433882 578898 433884 579134
rect 433644 578866 433884 578898
rect 439430 579454 439670 579486
rect 439430 579218 439432 579454
rect 439668 579218 439670 579454
rect 439430 579134 439670 579218
rect 439430 578898 439432 579134
rect 439668 578898 439670 579134
rect 439430 578866 439670 578898
rect 456608 579454 456848 579486
rect 456608 579218 456610 579454
rect 456846 579218 456848 579454
rect 456608 579134 456848 579218
rect 456608 578898 456610 579134
rect 456846 578898 456848 579134
rect 456608 578866 456848 578898
rect 477276 579454 477624 579486
rect 477276 579218 477332 579454
rect 477568 579218 477624 579454
rect 477276 579134 477624 579218
rect 477276 578898 477332 579134
rect 477568 578898 477624 579134
rect 477276 578866 477624 578898
rect 570980 579454 571328 579486
rect 570980 579218 571036 579454
rect 571272 579218 571328 579454
rect 570980 579134 571328 579218
rect 570980 578898 571036 579134
rect 571272 578898 571328 579134
rect 570980 578866 571328 578898
rect 578488 579454 579088 579486
rect 578488 579218 578670 579454
rect 578906 579218 579088 579454
rect 578488 579134 579088 579218
rect 578488 578898 578670 579134
rect 578906 578898 579088 579134
rect 578488 578866 579088 578898
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 4400 561454 5000 561486
rect 4400 561218 4582 561454
rect 4818 561218 5000 561454
rect 4400 561134 5000 561218
rect 4400 560898 4582 561134
rect 4818 560898 5000 561134
rect 4400 560866 5000 560898
rect 12296 561454 12644 561486
rect 12296 561218 12352 561454
rect 12588 561218 12644 561454
rect 12296 561134 12644 561218
rect 12296 560898 12352 561134
rect 12588 560898 12644 561134
rect 12296 560866 12644 560898
rect 107360 561454 107708 561486
rect 107360 561218 107416 561454
rect 107652 561218 107708 561454
rect 107360 561134 107708 561218
rect 107360 560898 107416 561134
rect 107652 560898 107708 561134
rect 107360 560866 107708 560898
rect 127056 561454 127296 561486
rect 127056 561218 127058 561454
rect 127294 561218 127296 561454
rect 127056 561134 127296 561218
rect 127056 560898 127058 561134
rect 127294 560898 127296 561134
rect 127056 560866 127296 560898
rect 140294 561454 140534 561486
rect 140294 561218 140296 561454
rect 140532 561218 140534 561454
rect 140294 561134 140534 561218
rect 140294 560898 140296 561134
rect 140532 560898 140534 561134
rect 140294 560866 140534 560898
rect 141100 561454 141340 561486
rect 141100 561218 141102 561454
rect 141338 561218 141340 561454
rect 141100 561134 141340 561218
rect 141100 560898 141102 561134
rect 141338 560898 141340 561134
rect 141100 560866 141340 560898
rect 147646 561454 147886 561486
rect 147646 561218 147648 561454
rect 147884 561218 147886 561454
rect 147646 561134 147886 561218
rect 147646 560898 147648 561134
rect 147884 560898 147886 561134
rect 147646 560866 147886 560898
rect 149298 561454 149538 561486
rect 149298 561218 149300 561454
rect 149536 561218 149538 561454
rect 149298 561134 149538 561218
rect 149298 560898 149300 561134
rect 149536 560898 149538 561134
rect 149298 560866 149538 560898
rect 150104 561454 150344 561486
rect 150104 561218 150106 561454
rect 150342 561218 150344 561454
rect 150104 561134 150344 561218
rect 150104 560898 150106 561134
rect 150342 560898 150344 561134
rect 150104 560866 150344 560898
rect 159104 561454 159344 561486
rect 159104 561218 159106 561454
rect 159342 561218 159344 561454
rect 159104 561134 159344 561218
rect 159104 560898 159106 561134
rect 159342 560898 159344 561134
rect 159104 560866 159344 560898
rect 168104 561454 168344 561486
rect 168104 561218 168106 561454
rect 168342 561218 168344 561454
rect 168104 561134 168344 561218
rect 168104 560898 168106 561134
rect 168342 560898 168344 561134
rect 168104 560866 168344 560898
rect 177104 561454 177344 561486
rect 177104 561218 177106 561454
rect 177342 561218 177344 561454
rect 177104 561134 177344 561218
rect 177104 560898 177106 561134
rect 177342 560898 177344 561134
rect 177104 560866 177344 560898
rect 186104 561454 186344 561486
rect 186104 561218 186106 561454
rect 186342 561218 186344 561454
rect 186104 561134 186344 561218
rect 186104 560898 186106 561134
rect 186342 560898 186344 561134
rect 186104 560866 186344 560898
rect 188666 561454 188906 561486
rect 188666 561218 188668 561454
rect 188904 561218 188906 561454
rect 188666 561134 188906 561218
rect 188666 560898 188668 561134
rect 188904 560898 188906 561134
rect 188666 560866 188906 560898
rect 190318 561454 190558 561486
rect 190318 561218 190320 561454
rect 190556 561218 190558 561454
rect 190318 561134 190558 561218
rect 190318 560898 190320 561134
rect 190556 560898 190558 561134
rect 190318 560866 190558 560898
rect 191124 561454 191364 561486
rect 191124 561218 191126 561454
rect 191362 561218 191364 561454
rect 191124 561134 191364 561218
rect 191124 560898 191126 561134
rect 191362 560898 191364 561134
rect 191124 560866 191364 560898
rect 200124 561454 200364 561486
rect 200124 561218 200126 561454
rect 200362 561218 200364 561454
rect 200124 561134 200364 561218
rect 200124 560898 200126 561134
rect 200362 560898 200364 561134
rect 200124 560866 200364 560898
rect 209124 561454 209364 561486
rect 209124 561218 209126 561454
rect 209362 561218 209364 561454
rect 209124 561134 209364 561218
rect 209124 560898 209126 561134
rect 209362 560898 209364 561134
rect 209124 560866 209364 560898
rect 218124 561454 218364 561486
rect 218124 561218 218126 561454
rect 218362 561218 218364 561454
rect 218124 561134 218364 561218
rect 218124 560898 218126 561134
rect 218362 560898 218364 561134
rect 218124 560866 218364 560898
rect 227124 561454 227364 561486
rect 227124 561218 227126 561454
rect 227362 561218 227364 561454
rect 227124 561134 227364 561218
rect 227124 560898 227126 561134
rect 227362 560898 227364 561134
rect 227124 560866 227364 560898
rect 229686 561454 229926 561486
rect 229686 561218 229688 561454
rect 229924 561218 229926 561454
rect 229686 561134 229926 561218
rect 229686 560898 229688 561134
rect 229924 560898 229926 561134
rect 229686 560866 229926 560898
rect 230338 561454 230578 561486
rect 230338 561218 230340 561454
rect 230576 561218 230578 561454
rect 230338 561134 230578 561218
rect 230338 560898 230340 561134
rect 230576 560898 230578 561134
rect 230338 560866 230578 560898
rect 231144 561454 231384 561486
rect 231144 561218 231146 561454
rect 231382 561218 231384 561454
rect 231144 561134 231384 561218
rect 231144 560898 231146 561134
rect 231382 560898 231384 561134
rect 231144 560866 231384 560898
rect 240144 561454 240384 561486
rect 240144 561218 240146 561454
rect 240382 561218 240384 561454
rect 240144 561134 240384 561218
rect 240144 560898 240146 561134
rect 240382 560898 240384 561134
rect 240144 560866 240384 560898
rect 249144 561454 249384 561486
rect 249144 561218 249146 561454
rect 249382 561218 249384 561454
rect 249144 561134 249384 561218
rect 249144 560898 249146 561134
rect 249382 560898 249384 561134
rect 249144 560866 249384 560898
rect 258144 561454 258384 561486
rect 258144 561218 258146 561454
rect 258382 561218 258384 561454
rect 258144 561134 258384 561218
rect 258144 560898 258146 561134
rect 258382 560898 258384 561134
rect 258144 560866 258384 560898
rect 267144 561454 267384 561486
rect 267144 561218 267146 561454
rect 267382 561218 267384 561454
rect 267144 561134 267384 561218
rect 267144 560898 267146 561134
rect 267382 560898 267384 561134
rect 267144 560866 267384 560898
rect 269706 561454 269946 561486
rect 269706 561218 269708 561454
rect 269944 561218 269946 561454
rect 269706 561134 269946 561218
rect 269706 560898 269708 561134
rect 269944 560898 269946 561134
rect 269706 560866 269946 560898
rect 270358 561454 270598 561486
rect 270358 561218 270360 561454
rect 270596 561218 270598 561454
rect 270358 561134 270598 561218
rect 270358 560898 270360 561134
rect 270596 560898 270598 561134
rect 270358 560866 270598 560898
rect 271164 561454 271404 561486
rect 271164 561218 271166 561454
rect 271402 561218 271404 561454
rect 271164 561134 271404 561218
rect 271164 560898 271166 561134
rect 271402 560898 271404 561134
rect 271164 560866 271404 560898
rect 280164 561454 280404 561486
rect 280164 561218 280166 561454
rect 280402 561218 280404 561454
rect 280164 561134 280404 561218
rect 280164 560898 280166 561134
rect 280402 560898 280404 561134
rect 280164 560866 280404 560898
rect 289164 561454 289404 561486
rect 289164 561218 289166 561454
rect 289402 561218 289404 561454
rect 289164 561134 289404 561218
rect 289164 560898 289166 561134
rect 289402 560898 289404 561134
rect 289164 560866 289404 560898
rect 298164 561454 298404 561486
rect 298164 561218 298166 561454
rect 298402 561218 298404 561454
rect 298164 561134 298404 561218
rect 298164 560898 298166 561134
rect 298402 560898 298404 561134
rect 298164 560866 298404 560898
rect 307164 561454 307404 561486
rect 307164 561218 307166 561454
rect 307402 561218 307404 561454
rect 307164 561134 307404 561218
rect 307164 560898 307166 561134
rect 307402 560898 307404 561134
rect 307164 560866 307404 560898
rect 309726 561454 309966 561486
rect 309726 561218 309728 561454
rect 309964 561218 309966 561454
rect 309726 561134 309966 561218
rect 309726 560898 309728 561134
rect 309964 560898 309966 561134
rect 309726 560866 309966 560898
rect 311378 561454 311618 561486
rect 311378 561218 311380 561454
rect 311616 561218 311618 561454
rect 311378 561134 311618 561218
rect 311378 560898 311380 561134
rect 311616 560898 311618 561134
rect 311378 560866 311618 560898
rect 312184 561454 312424 561486
rect 312184 561218 312186 561454
rect 312422 561218 312424 561454
rect 312184 561134 312424 561218
rect 312184 560898 312186 561134
rect 312422 560898 312424 561134
rect 312184 560866 312424 560898
rect 321184 561454 321424 561486
rect 321184 561218 321186 561454
rect 321422 561218 321424 561454
rect 321184 561134 321424 561218
rect 321184 560898 321186 561134
rect 321422 560898 321424 561134
rect 321184 560866 321424 560898
rect 330184 561454 330424 561486
rect 330184 561218 330186 561454
rect 330422 561218 330424 561454
rect 330184 561134 330424 561218
rect 330184 560898 330186 561134
rect 330422 560898 330424 561134
rect 330184 560866 330424 560898
rect 339184 561454 339424 561486
rect 339184 561218 339186 561454
rect 339422 561218 339424 561454
rect 339184 561134 339424 561218
rect 339184 560898 339186 561134
rect 339422 560898 339424 561134
rect 339184 560866 339424 560898
rect 348184 561454 348424 561486
rect 348184 561218 348186 561454
rect 348422 561218 348424 561454
rect 348184 561134 348424 561218
rect 348184 560898 348186 561134
rect 348422 560898 348424 561134
rect 348184 560866 348424 560898
rect 350746 561454 350986 561486
rect 350746 561218 350748 561454
rect 350984 561218 350986 561454
rect 350746 561134 350986 561218
rect 350746 560898 350748 561134
rect 350984 560898 350986 561134
rect 350746 560866 350986 560898
rect 352398 561454 352638 561486
rect 352398 561218 352400 561454
rect 352636 561218 352638 561454
rect 352398 561134 352638 561218
rect 352398 560898 352400 561134
rect 352636 560898 352638 561134
rect 352398 560866 352638 560898
rect 353204 561454 353444 561486
rect 353204 561218 353206 561454
rect 353442 561218 353444 561454
rect 353204 561134 353444 561218
rect 353204 560898 353206 561134
rect 353442 560898 353444 561134
rect 353204 560866 353444 560898
rect 362204 561454 362444 561486
rect 362204 561218 362206 561454
rect 362442 561218 362444 561454
rect 362204 561134 362444 561218
rect 362204 560898 362206 561134
rect 362442 560898 362444 561134
rect 362204 560866 362444 560898
rect 371204 561454 371444 561486
rect 371204 561218 371206 561454
rect 371442 561218 371444 561454
rect 371204 561134 371444 561218
rect 371204 560898 371206 561134
rect 371442 560898 371444 561134
rect 371204 560866 371444 560898
rect 380204 561454 380444 561486
rect 380204 561218 380206 561454
rect 380442 561218 380444 561454
rect 380204 561134 380444 561218
rect 380204 560898 380206 561134
rect 380442 560898 380444 561134
rect 380204 560866 380444 560898
rect 389204 561454 389444 561486
rect 389204 561218 389206 561454
rect 389442 561218 389444 561454
rect 389204 561134 389444 561218
rect 389204 560898 389206 561134
rect 389442 560898 389444 561134
rect 389204 560866 389444 560898
rect 391766 561454 392006 561486
rect 391766 561218 391768 561454
rect 392004 561218 392006 561454
rect 391766 561134 392006 561218
rect 391766 560898 391768 561134
rect 392004 560898 392006 561134
rect 391766 560866 392006 560898
rect 392418 561454 392658 561486
rect 392418 561218 392420 561454
rect 392656 561218 392658 561454
rect 392418 561134 392658 561218
rect 392418 560898 392420 561134
rect 392656 560898 392658 561134
rect 392418 560866 392658 560898
rect 393224 561454 393464 561486
rect 393224 561218 393226 561454
rect 393462 561218 393464 561454
rect 393224 561134 393464 561218
rect 393224 560898 393226 561134
rect 393462 560898 393464 561134
rect 393224 560866 393464 560898
rect 402224 561454 402464 561486
rect 402224 561218 402226 561454
rect 402462 561218 402464 561454
rect 402224 561134 402464 561218
rect 402224 560898 402226 561134
rect 402462 560898 402464 561134
rect 402224 560866 402464 560898
rect 411224 561454 411464 561486
rect 411224 561218 411226 561454
rect 411462 561218 411464 561454
rect 411224 561134 411464 561218
rect 411224 560898 411226 561134
rect 411462 560898 411464 561134
rect 411224 560866 411464 560898
rect 420224 561454 420464 561486
rect 420224 561218 420226 561454
rect 420462 561218 420464 561454
rect 420224 561134 420464 561218
rect 420224 560898 420226 561134
rect 420462 560898 420464 561134
rect 420224 560866 420464 560898
rect 429224 561454 429464 561486
rect 429224 561218 429226 561454
rect 429462 561218 429464 561454
rect 429224 561134 429464 561218
rect 429224 560898 429226 561134
rect 429462 560898 429464 561134
rect 429224 560866 429464 560898
rect 431786 561454 432026 561486
rect 431786 561218 431788 561454
rect 432024 561218 432026 561454
rect 431786 561134 432026 561218
rect 431786 560898 431788 561134
rect 432024 560898 432026 561134
rect 431786 560866 432026 560898
rect 432438 561454 432678 561486
rect 432438 561218 432440 561454
rect 432676 561218 432678 561454
rect 432438 561134 432678 561218
rect 432438 560898 432440 561134
rect 432676 560898 432678 561134
rect 432438 560866 432678 560898
rect 433244 561454 433484 561486
rect 433244 561218 433246 561454
rect 433482 561218 433484 561454
rect 433244 561134 433484 561218
rect 433244 560898 433246 561134
rect 433482 560898 433484 561134
rect 433244 560866 433484 560898
rect 439790 561454 440030 561486
rect 439790 561218 439792 561454
rect 440028 561218 440030 561454
rect 439790 561134 440030 561218
rect 439790 560898 439792 561134
rect 440028 560898 440030 561134
rect 439790 560866 440030 560898
rect 457008 561454 457248 561486
rect 457008 561218 457010 561454
rect 457246 561218 457248 561454
rect 457008 561134 457248 561218
rect 457008 560898 457010 561134
rect 457246 560898 457248 561134
rect 457008 560866 457248 560898
rect 476596 561454 476944 561486
rect 476596 561218 476652 561454
rect 476888 561218 476944 561454
rect 476596 561134 476944 561218
rect 476596 560898 476652 561134
rect 476888 560898 476944 561134
rect 476596 560866 476944 560898
rect 571660 561454 572008 561486
rect 571660 561218 571716 561454
rect 571952 561218 572008 561454
rect 571660 561134 572008 561218
rect 571660 560898 571716 561134
rect 571952 560898 572008 561134
rect 571660 560866 572008 560898
rect 579288 561454 579888 561486
rect 579288 561218 579470 561454
rect 579706 561218 579888 561454
rect 579288 561134 579888 561218
rect 579288 560898 579470 561134
rect 579706 560898 579888 561134
rect 579288 560866 579888 560898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect 5200 543454 5800 543486
rect 5200 543218 5382 543454
rect 5618 543218 5800 543454
rect 5200 543134 5800 543218
rect 5200 542898 5382 543134
rect 5618 542898 5800 543134
rect 5200 542866 5800 542898
rect 127456 543454 127696 543486
rect 127456 543218 127458 543454
rect 127694 543218 127696 543454
rect 127456 543134 127696 543218
rect 127456 542898 127458 543134
rect 127694 542898 127696 543134
rect 127456 542866 127696 542898
rect 140654 543454 140894 543486
rect 140654 543218 140656 543454
rect 140892 543218 140894 543454
rect 140654 543134 140894 543218
rect 140654 542898 140656 543134
rect 140892 542898 140894 543134
rect 140654 542866 140894 542898
rect 141500 543454 141740 543486
rect 141500 543218 141502 543454
rect 141738 543218 141740 543454
rect 141500 543134 141740 543218
rect 141500 542898 141502 543134
rect 141738 542898 141740 543134
rect 141500 542866 141740 542898
rect 147286 543454 147526 543486
rect 147286 543218 147288 543454
rect 147524 543218 147526 543454
rect 147286 543134 147526 543218
rect 147286 542898 147288 543134
rect 147524 542898 147526 543134
rect 147286 542866 147526 542898
rect 149658 543454 149898 543486
rect 149658 543218 149660 543454
rect 149896 543218 149898 543454
rect 149658 543134 149898 543218
rect 149658 542898 149660 543134
rect 149896 542898 149898 543134
rect 149658 542866 149898 542898
rect 150504 543454 150744 543486
rect 150504 543218 150506 543454
rect 150742 543218 150744 543454
rect 150504 543134 150744 543218
rect 150504 542898 150506 543134
rect 150742 542898 150744 543134
rect 150504 542866 150744 542898
rect 159504 543454 159744 543486
rect 159504 543218 159506 543454
rect 159742 543218 159744 543454
rect 159504 543134 159744 543218
rect 159504 542898 159506 543134
rect 159742 542898 159744 543134
rect 159504 542866 159744 542898
rect 168504 543454 168744 543486
rect 168504 543218 168506 543454
rect 168742 543218 168744 543454
rect 168504 543134 168744 543218
rect 168504 542898 168506 543134
rect 168742 542898 168744 543134
rect 168504 542866 168744 542898
rect 177504 543454 177744 543486
rect 177504 543218 177506 543454
rect 177742 543218 177744 543454
rect 177504 543134 177744 543218
rect 177504 542898 177506 543134
rect 177742 542898 177744 543134
rect 177504 542866 177744 542898
rect 186504 543454 186744 543486
rect 186504 543218 186506 543454
rect 186742 543218 186744 543454
rect 186504 543134 186744 543218
rect 186504 542898 186506 543134
rect 186742 542898 186744 543134
rect 186504 542866 186744 542898
rect 188306 543454 188546 543486
rect 188306 543218 188308 543454
rect 188544 543218 188546 543454
rect 188306 543134 188546 543218
rect 188306 542898 188308 543134
rect 188544 542898 188546 543134
rect 188306 542866 188546 542898
rect 190678 543454 190918 543486
rect 190678 543218 190680 543454
rect 190916 543218 190918 543454
rect 190678 543134 190918 543218
rect 190678 542898 190680 543134
rect 190916 542898 190918 543134
rect 190678 542866 190918 542898
rect 191524 543454 191764 543486
rect 191524 543218 191526 543454
rect 191762 543218 191764 543454
rect 191524 543134 191764 543218
rect 191524 542898 191526 543134
rect 191762 542898 191764 543134
rect 191524 542866 191764 542898
rect 200524 543454 200764 543486
rect 200524 543218 200526 543454
rect 200762 543218 200764 543454
rect 200524 543134 200764 543218
rect 200524 542898 200526 543134
rect 200762 542898 200764 543134
rect 200524 542866 200764 542898
rect 209524 543454 209764 543486
rect 209524 543218 209526 543454
rect 209762 543218 209764 543454
rect 209524 543134 209764 543218
rect 209524 542898 209526 543134
rect 209762 542898 209764 543134
rect 209524 542866 209764 542898
rect 218524 543454 218764 543486
rect 218524 543218 218526 543454
rect 218762 543218 218764 543454
rect 218524 543134 218764 543218
rect 218524 542898 218526 543134
rect 218762 542898 218764 543134
rect 218524 542866 218764 542898
rect 227524 543454 227764 543486
rect 227524 543218 227526 543454
rect 227762 543218 227764 543454
rect 227524 543134 227764 543218
rect 227524 542898 227526 543134
rect 227762 542898 227764 543134
rect 227524 542866 227764 542898
rect 229326 543454 229566 543486
rect 229326 543218 229328 543454
rect 229564 543218 229566 543454
rect 229326 543134 229566 543218
rect 229326 542898 229328 543134
rect 229564 542898 229566 543134
rect 229326 542866 229566 542898
rect 230698 543454 230938 543486
rect 230698 543218 230700 543454
rect 230936 543218 230938 543454
rect 230698 543134 230938 543218
rect 230698 542898 230700 543134
rect 230936 542898 230938 543134
rect 230698 542866 230938 542898
rect 231544 543454 231784 543486
rect 231544 543218 231546 543454
rect 231782 543218 231784 543454
rect 231544 543134 231784 543218
rect 231544 542898 231546 543134
rect 231782 542898 231784 543134
rect 231544 542866 231784 542898
rect 240544 543454 240784 543486
rect 240544 543218 240546 543454
rect 240782 543218 240784 543454
rect 240544 543134 240784 543218
rect 240544 542898 240546 543134
rect 240782 542898 240784 543134
rect 240544 542866 240784 542898
rect 249544 543454 249784 543486
rect 249544 543218 249546 543454
rect 249782 543218 249784 543454
rect 249544 543134 249784 543218
rect 249544 542898 249546 543134
rect 249782 542898 249784 543134
rect 249544 542866 249784 542898
rect 258544 543454 258784 543486
rect 258544 543218 258546 543454
rect 258782 543218 258784 543454
rect 258544 543134 258784 543218
rect 258544 542898 258546 543134
rect 258782 542898 258784 543134
rect 258544 542866 258784 542898
rect 267544 543454 267784 543486
rect 267544 543218 267546 543454
rect 267782 543218 267784 543454
rect 267544 543134 267784 543218
rect 267544 542898 267546 543134
rect 267782 542898 267784 543134
rect 267544 542866 267784 542898
rect 269346 543454 269586 543486
rect 269346 543218 269348 543454
rect 269584 543218 269586 543454
rect 269346 543134 269586 543218
rect 269346 542898 269348 543134
rect 269584 542898 269586 543134
rect 269346 542866 269586 542898
rect 270718 543454 270958 543486
rect 270718 543218 270720 543454
rect 270956 543218 270958 543454
rect 270718 543134 270958 543218
rect 270718 542898 270720 543134
rect 270956 542898 270958 543134
rect 270718 542866 270958 542898
rect 271564 543454 271804 543486
rect 271564 543218 271566 543454
rect 271802 543218 271804 543454
rect 271564 543134 271804 543218
rect 271564 542898 271566 543134
rect 271802 542898 271804 543134
rect 271564 542866 271804 542898
rect 280564 543454 280804 543486
rect 280564 543218 280566 543454
rect 280802 543218 280804 543454
rect 280564 543134 280804 543218
rect 280564 542898 280566 543134
rect 280802 542898 280804 543134
rect 280564 542866 280804 542898
rect 289564 543454 289804 543486
rect 289564 543218 289566 543454
rect 289802 543218 289804 543454
rect 289564 543134 289804 543218
rect 289564 542898 289566 543134
rect 289802 542898 289804 543134
rect 289564 542866 289804 542898
rect 298564 543454 298804 543486
rect 298564 543218 298566 543454
rect 298802 543218 298804 543454
rect 298564 543134 298804 543218
rect 298564 542898 298566 543134
rect 298802 542898 298804 543134
rect 298564 542866 298804 542898
rect 307564 543454 307804 543486
rect 307564 543218 307566 543454
rect 307802 543218 307804 543454
rect 307564 543134 307804 543218
rect 307564 542898 307566 543134
rect 307802 542898 307804 543134
rect 307564 542866 307804 542898
rect 309366 543454 309606 543486
rect 309366 543218 309368 543454
rect 309604 543218 309606 543454
rect 309366 543134 309606 543218
rect 309366 542898 309368 543134
rect 309604 542898 309606 543134
rect 309366 542866 309606 542898
rect 311738 543454 311978 543486
rect 311738 543218 311740 543454
rect 311976 543218 311978 543454
rect 311738 543134 311978 543218
rect 311738 542898 311740 543134
rect 311976 542898 311978 543134
rect 311738 542866 311978 542898
rect 312584 543454 312824 543486
rect 312584 543218 312586 543454
rect 312822 543218 312824 543454
rect 312584 543134 312824 543218
rect 312584 542898 312586 543134
rect 312822 542898 312824 543134
rect 312584 542866 312824 542898
rect 321584 543454 321824 543486
rect 321584 543218 321586 543454
rect 321822 543218 321824 543454
rect 321584 543134 321824 543218
rect 321584 542898 321586 543134
rect 321822 542898 321824 543134
rect 321584 542866 321824 542898
rect 330584 543454 330824 543486
rect 330584 543218 330586 543454
rect 330822 543218 330824 543454
rect 330584 543134 330824 543218
rect 330584 542898 330586 543134
rect 330822 542898 330824 543134
rect 330584 542866 330824 542898
rect 339584 543454 339824 543486
rect 339584 543218 339586 543454
rect 339822 543218 339824 543454
rect 339584 543134 339824 543218
rect 339584 542898 339586 543134
rect 339822 542898 339824 543134
rect 339584 542866 339824 542898
rect 348584 543454 348824 543486
rect 348584 543218 348586 543454
rect 348822 543218 348824 543454
rect 348584 543134 348824 543218
rect 348584 542898 348586 543134
rect 348822 542898 348824 543134
rect 348584 542866 348824 542898
rect 350386 543454 350626 543486
rect 350386 543218 350388 543454
rect 350624 543218 350626 543454
rect 350386 543134 350626 543218
rect 350386 542898 350388 543134
rect 350624 542898 350626 543134
rect 350386 542866 350626 542898
rect 352758 543454 352998 543486
rect 352758 543218 352760 543454
rect 352996 543218 352998 543454
rect 352758 543134 352998 543218
rect 352758 542898 352760 543134
rect 352996 542898 352998 543134
rect 352758 542866 352998 542898
rect 353604 543454 353844 543486
rect 353604 543218 353606 543454
rect 353842 543218 353844 543454
rect 353604 543134 353844 543218
rect 353604 542898 353606 543134
rect 353842 542898 353844 543134
rect 353604 542866 353844 542898
rect 362604 543454 362844 543486
rect 362604 543218 362606 543454
rect 362842 543218 362844 543454
rect 362604 543134 362844 543218
rect 362604 542898 362606 543134
rect 362842 542898 362844 543134
rect 362604 542866 362844 542898
rect 371604 543454 371844 543486
rect 371604 543218 371606 543454
rect 371842 543218 371844 543454
rect 371604 543134 371844 543218
rect 371604 542898 371606 543134
rect 371842 542898 371844 543134
rect 371604 542866 371844 542898
rect 380604 543454 380844 543486
rect 380604 543218 380606 543454
rect 380842 543218 380844 543454
rect 380604 543134 380844 543218
rect 380604 542898 380606 543134
rect 380842 542898 380844 543134
rect 380604 542866 380844 542898
rect 389604 543454 389844 543486
rect 389604 543218 389606 543454
rect 389842 543218 389844 543454
rect 389604 543134 389844 543218
rect 389604 542898 389606 543134
rect 389842 542898 389844 543134
rect 389604 542866 389844 542898
rect 391406 543454 391646 543486
rect 391406 543218 391408 543454
rect 391644 543218 391646 543454
rect 391406 543134 391646 543218
rect 391406 542898 391408 543134
rect 391644 542898 391646 543134
rect 391406 542866 391646 542898
rect 392778 543454 393018 543486
rect 392778 543218 392780 543454
rect 393016 543218 393018 543454
rect 392778 543134 393018 543218
rect 392778 542898 392780 543134
rect 393016 542898 393018 543134
rect 392778 542866 393018 542898
rect 393624 543454 393864 543486
rect 393624 543218 393626 543454
rect 393862 543218 393864 543454
rect 393624 543134 393864 543218
rect 393624 542898 393626 543134
rect 393862 542898 393864 543134
rect 393624 542866 393864 542898
rect 402624 543454 402864 543486
rect 402624 543218 402626 543454
rect 402862 543218 402864 543454
rect 402624 543134 402864 543218
rect 402624 542898 402626 543134
rect 402862 542898 402864 543134
rect 402624 542866 402864 542898
rect 411624 543454 411864 543486
rect 411624 543218 411626 543454
rect 411862 543218 411864 543454
rect 411624 543134 411864 543218
rect 411624 542898 411626 543134
rect 411862 542898 411864 543134
rect 411624 542866 411864 542898
rect 420624 543454 420864 543486
rect 420624 543218 420626 543454
rect 420862 543218 420864 543454
rect 420624 543134 420864 543218
rect 420624 542898 420626 543134
rect 420862 542898 420864 543134
rect 420624 542866 420864 542898
rect 429624 543454 429864 543486
rect 429624 543218 429626 543454
rect 429862 543218 429864 543454
rect 429624 543134 429864 543218
rect 429624 542898 429626 543134
rect 429862 542898 429864 543134
rect 429624 542866 429864 542898
rect 431426 543454 431666 543486
rect 431426 543218 431428 543454
rect 431664 543218 431666 543454
rect 431426 543134 431666 543218
rect 431426 542898 431428 543134
rect 431664 542898 431666 543134
rect 431426 542866 431666 542898
rect 432798 543454 433038 543486
rect 432798 543218 432800 543454
rect 433036 543218 433038 543454
rect 432798 543134 433038 543218
rect 432798 542898 432800 543134
rect 433036 542898 433038 543134
rect 432798 542866 433038 542898
rect 433644 543454 433884 543486
rect 433644 543218 433646 543454
rect 433882 543218 433884 543454
rect 433644 543134 433884 543218
rect 433644 542898 433646 543134
rect 433882 542898 433884 543134
rect 433644 542866 433884 542898
rect 439430 543454 439670 543486
rect 439430 543218 439432 543454
rect 439668 543218 439670 543454
rect 439430 543134 439670 543218
rect 439430 542898 439432 543134
rect 439668 542898 439670 543134
rect 439430 542866 439670 542898
rect 456608 543454 456848 543486
rect 456608 543218 456610 543454
rect 456846 543218 456848 543454
rect 456608 543134 456848 543218
rect 456608 542898 456610 543134
rect 456846 542898 456848 543134
rect 456608 542866 456848 542898
rect 578488 543454 579088 543486
rect 578488 543218 578670 543454
rect 578906 543218 579088 543454
rect 578488 543134 579088 543218
rect 578488 542898 578670 543134
rect 578906 542898 579088 543134
rect 578488 542866 579088 542898
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 4400 525454 5000 525486
rect 4400 525218 4582 525454
rect 4818 525218 5000 525454
rect 4400 525134 5000 525218
rect 4400 524898 4582 525134
rect 4818 524898 5000 525134
rect 4400 524866 5000 524898
rect 127056 525454 127296 525486
rect 127056 525218 127058 525454
rect 127294 525218 127296 525454
rect 127056 525134 127296 525218
rect 127056 524898 127058 525134
rect 127294 524898 127296 525134
rect 127056 524866 127296 524898
rect 140294 525454 140534 525486
rect 140294 525218 140296 525454
rect 140532 525218 140534 525454
rect 140294 525134 140534 525218
rect 140294 524898 140296 525134
rect 140532 524898 140534 525134
rect 140294 524866 140534 524898
rect 141100 525454 141340 525486
rect 141100 525218 141102 525454
rect 141338 525218 141340 525454
rect 141100 525134 141340 525218
rect 141100 524898 141102 525134
rect 141338 524898 141340 525134
rect 141100 524866 141340 524898
rect 147646 525454 147886 525486
rect 147646 525218 147648 525454
rect 147884 525218 147886 525454
rect 147646 525134 147886 525218
rect 147646 524898 147648 525134
rect 147884 524898 147886 525134
rect 147646 524866 147886 524898
rect 149298 525454 149538 525486
rect 149298 525218 149300 525454
rect 149536 525218 149538 525454
rect 149298 525134 149538 525218
rect 149298 524898 149300 525134
rect 149536 524898 149538 525134
rect 149298 524866 149538 524898
rect 150104 525454 150344 525486
rect 150104 525218 150106 525454
rect 150342 525218 150344 525454
rect 150104 525134 150344 525218
rect 150104 524898 150106 525134
rect 150342 524898 150344 525134
rect 150104 524866 150344 524898
rect 159104 525454 159344 525486
rect 159104 525218 159106 525454
rect 159342 525218 159344 525454
rect 159104 525134 159344 525218
rect 159104 524898 159106 525134
rect 159342 524898 159344 525134
rect 159104 524866 159344 524898
rect 168104 525454 168344 525486
rect 168104 525218 168106 525454
rect 168342 525218 168344 525454
rect 168104 525134 168344 525218
rect 168104 524898 168106 525134
rect 168342 524898 168344 525134
rect 168104 524866 168344 524898
rect 177104 525454 177344 525486
rect 177104 525218 177106 525454
rect 177342 525218 177344 525454
rect 177104 525134 177344 525218
rect 177104 524898 177106 525134
rect 177342 524898 177344 525134
rect 177104 524866 177344 524898
rect 186104 525454 186344 525486
rect 186104 525218 186106 525454
rect 186342 525218 186344 525454
rect 186104 525134 186344 525218
rect 186104 524898 186106 525134
rect 186342 524898 186344 525134
rect 186104 524866 186344 524898
rect 188666 525454 188906 525486
rect 188666 525218 188668 525454
rect 188904 525218 188906 525454
rect 188666 525134 188906 525218
rect 188666 524898 188668 525134
rect 188904 524898 188906 525134
rect 188666 524866 188906 524898
rect 190318 525454 190558 525486
rect 190318 525218 190320 525454
rect 190556 525218 190558 525454
rect 190318 525134 190558 525218
rect 190318 524898 190320 525134
rect 190556 524898 190558 525134
rect 190318 524866 190558 524898
rect 191124 525454 191364 525486
rect 191124 525218 191126 525454
rect 191362 525218 191364 525454
rect 191124 525134 191364 525218
rect 191124 524898 191126 525134
rect 191362 524898 191364 525134
rect 191124 524866 191364 524898
rect 200124 525454 200364 525486
rect 200124 525218 200126 525454
rect 200362 525218 200364 525454
rect 200124 525134 200364 525218
rect 200124 524898 200126 525134
rect 200362 524898 200364 525134
rect 200124 524866 200364 524898
rect 209124 525454 209364 525486
rect 209124 525218 209126 525454
rect 209362 525218 209364 525454
rect 209124 525134 209364 525218
rect 209124 524898 209126 525134
rect 209362 524898 209364 525134
rect 209124 524866 209364 524898
rect 218124 525454 218364 525486
rect 218124 525218 218126 525454
rect 218362 525218 218364 525454
rect 218124 525134 218364 525218
rect 218124 524898 218126 525134
rect 218362 524898 218364 525134
rect 218124 524866 218364 524898
rect 227124 525454 227364 525486
rect 227124 525218 227126 525454
rect 227362 525218 227364 525454
rect 227124 525134 227364 525218
rect 227124 524898 227126 525134
rect 227362 524898 227364 525134
rect 227124 524866 227364 524898
rect 229686 525454 229926 525486
rect 229686 525218 229688 525454
rect 229924 525218 229926 525454
rect 229686 525134 229926 525218
rect 229686 524898 229688 525134
rect 229924 524898 229926 525134
rect 229686 524866 229926 524898
rect 230338 525454 230578 525486
rect 230338 525218 230340 525454
rect 230576 525218 230578 525454
rect 230338 525134 230578 525218
rect 230338 524898 230340 525134
rect 230576 524898 230578 525134
rect 230338 524866 230578 524898
rect 231144 525454 231384 525486
rect 231144 525218 231146 525454
rect 231382 525218 231384 525454
rect 231144 525134 231384 525218
rect 231144 524898 231146 525134
rect 231382 524898 231384 525134
rect 231144 524866 231384 524898
rect 240144 525454 240384 525486
rect 240144 525218 240146 525454
rect 240382 525218 240384 525454
rect 240144 525134 240384 525218
rect 240144 524898 240146 525134
rect 240382 524898 240384 525134
rect 240144 524866 240384 524898
rect 249144 525454 249384 525486
rect 249144 525218 249146 525454
rect 249382 525218 249384 525454
rect 249144 525134 249384 525218
rect 249144 524898 249146 525134
rect 249382 524898 249384 525134
rect 249144 524866 249384 524898
rect 258144 525454 258384 525486
rect 258144 525218 258146 525454
rect 258382 525218 258384 525454
rect 258144 525134 258384 525218
rect 258144 524898 258146 525134
rect 258382 524898 258384 525134
rect 258144 524866 258384 524898
rect 267144 525454 267384 525486
rect 267144 525218 267146 525454
rect 267382 525218 267384 525454
rect 267144 525134 267384 525218
rect 267144 524898 267146 525134
rect 267382 524898 267384 525134
rect 267144 524866 267384 524898
rect 269706 525454 269946 525486
rect 269706 525218 269708 525454
rect 269944 525218 269946 525454
rect 269706 525134 269946 525218
rect 269706 524898 269708 525134
rect 269944 524898 269946 525134
rect 269706 524866 269946 524898
rect 270358 525454 270598 525486
rect 270358 525218 270360 525454
rect 270596 525218 270598 525454
rect 270358 525134 270598 525218
rect 270358 524898 270360 525134
rect 270596 524898 270598 525134
rect 270358 524866 270598 524898
rect 271164 525454 271404 525486
rect 271164 525218 271166 525454
rect 271402 525218 271404 525454
rect 271164 525134 271404 525218
rect 271164 524898 271166 525134
rect 271402 524898 271404 525134
rect 271164 524866 271404 524898
rect 280164 525454 280404 525486
rect 280164 525218 280166 525454
rect 280402 525218 280404 525454
rect 280164 525134 280404 525218
rect 280164 524898 280166 525134
rect 280402 524898 280404 525134
rect 280164 524866 280404 524898
rect 289164 525454 289404 525486
rect 289164 525218 289166 525454
rect 289402 525218 289404 525454
rect 289164 525134 289404 525218
rect 289164 524898 289166 525134
rect 289402 524898 289404 525134
rect 289164 524866 289404 524898
rect 298164 525454 298404 525486
rect 298164 525218 298166 525454
rect 298402 525218 298404 525454
rect 298164 525134 298404 525218
rect 298164 524898 298166 525134
rect 298402 524898 298404 525134
rect 298164 524866 298404 524898
rect 307164 525454 307404 525486
rect 307164 525218 307166 525454
rect 307402 525218 307404 525454
rect 307164 525134 307404 525218
rect 307164 524898 307166 525134
rect 307402 524898 307404 525134
rect 307164 524866 307404 524898
rect 309726 525454 309966 525486
rect 309726 525218 309728 525454
rect 309964 525218 309966 525454
rect 309726 525134 309966 525218
rect 309726 524898 309728 525134
rect 309964 524898 309966 525134
rect 309726 524866 309966 524898
rect 311378 525454 311618 525486
rect 311378 525218 311380 525454
rect 311616 525218 311618 525454
rect 311378 525134 311618 525218
rect 311378 524898 311380 525134
rect 311616 524898 311618 525134
rect 311378 524866 311618 524898
rect 312184 525454 312424 525486
rect 312184 525218 312186 525454
rect 312422 525218 312424 525454
rect 312184 525134 312424 525218
rect 312184 524898 312186 525134
rect 312422 524898 312424 525134
rect 312184 524866 312424 524898
rect 321184 525454 321424 525486
rect 321184 525218 321186 525454
rect 321422 525218 321424 525454
rect 321184 525134 321424 525218
rect 321184 524898 321186 525134
rect 321422 524898 321424 525134
rect 321184 524866 321424 524898
rect 330184 525454 330424 525486
rect 330184 525218 330186 525454
rect 330422 525218 330424 525454
rect 330184 525134 330424 525218
rect 330184 524898 330186 525134
rect 330422 524898 330424 525134
rect 330184 524866 330424 524898
rect 339184 525454 339424 525486
rect 339184 525218 339186 525454
rect 339422 525218 339424 525454
rect 339184 525134 339424 525218
rect 339184 524898 339186 525134
rect 339422 524898 339424 525134
rect 339184 524866 339424 524898
rect 348184 525454 348424 525486
rect 348184 525218 348186 525454
rect 348422 525218 348424 525454
rect 348184 525134 348424 525218
rect 348184 524898 348186 525134
rect 348422 524898 348424 525134
rect 348184 524866 348424 524898
rect 350746 525454 350986 525486
rect 350746 525218 350748 525454
rect 350984 525218 350986 525454
rect 350746 525134 350986 525218
rect 350746 524898 350748 525134
rect 350984 524898 350986 525134
rect 350746 524866 350986 524898
rect 352398 525454 352638 525486
rect 352398 525218 352400 525454
rect 352636 525218 352638 525454
rect 352398 525134 352638 525218
rect 352398 524898 352400 525134
rect 352636 524898 352638 525134
rect 352398 524866 352638 524898
rect 353204 525454 353444 525486
rect 353204 525218 353206 525454
rect 353442 525218 353444 525454
rect 353204 525134 353444 525218
rect 353204 524898 353206 525134
rect 353442 524898 353444 525134
rect 353204 524866 353444 524898
rect 362204 525454 362444 525486
rect 362204 525218 362206 525454
rect 362442 525218 362444 525454
rect 362204 525134 362444 525218
rect 362204 524898 362206 525134
rect 362442 524898 362444 525134
rect 362204 524866 362444 524898
rect 371204 525454 371444 525486
rect 371204 525218 371206 525454
rect 371442 525218 371444 525454
rect 371204 525134 371444 525218
rect 371204 524898 371206 525134
rect 371442 524898 371444 525134
rect 371204 524866 371444 524898
rect 380204 525454 380444 525486
rect 380204 525218 380206 525454
rect 380442 525218 380444 525454
rect 380204 525134 380444 525218
rect 380204 524898 380206 525134
rect 380442 524898 380444 525134
rect 380204 524866 380444 524898
rect 389204 525454 389444 525486
rect 389204 525218 389206 525454
rect 389442 525218 389444 525454
rect 389204 525134 389444 525218
rect 389204 524898 389206 525134
rect 389442 524898 389444 525134
rect 389204 524866 389444 524898
rect 391766 525454 392006 525486
rect 391766 525218 391768 525454
rect 392004 525218 392006 525454
rect 391766 525134 392006 525218
rect 391766 524898 391768 525134
rect 392004 524898 392006 525134
rect 391766 524866 392006 524898
rect 392418 525454 392658 525486
rect 392418 525218 392420 525454
rect 392656 525218 392658 525454
rect 392418 525134 392658 525218
rect 392418 524898 392420 525134
rect 392656 524898 392658 525134
rect 392418 524866 392658 524898
rect 393224 525454 393464 525486
rect 393224 525218 393226 525454
rect 393462 525218 393464 525454
rect 393224 525134 393464 525218
rect 393224 524898 393226 525134
rect 393462 524898 393464 525134
rect 393224 524866 393464 524898
rect 402224 525454 402464 525486
rect 402224 525218 402226 525454
rect 402462 525218 402464 525454
rect 402224 525134 402464 525218
rect 402224 524898 402226 525134
rect 402462 524898 402464 525134
rect 402224 524866 402464 524898
rect 411224 525454 411464 525486
rect 411224 525218 411226 525454
rect 411462 525218 411464 525454
rect 411224 525134 411464 525218
rect 411224 524898 411226 525134
rect 411462 524898 411464 525134
rect 411224 524866 411464 524898
rect 420224 525454 420464 525486
rect 420224 525218 420226 525454
rect 420462 525218 420464 525454
rect 420224 525134 420464 525218
rect 420224 524898 420226 525134
rect 420462 524898 420464 525134
rect 420224 524866 420464 524898
rect 429224 525454 429464 525486
rect 429224 525218 429226 525454
rect 429462 525218 429464 525454
rect 429224 525134 429464 525218
rect 429224 524898 429226 525134
rect 429462 524898 429464 525134
rect 429224 524866 429464 524898
rect 431786 525454 432026 525486
rect 431786 525218 431788 525454
rect 432024 525218 432026 525454
rect 431786 525134 432026 525218
rect 431786 524898 431788 525134
rect 432024 524898 432026 525134
rect 431786 524866 432026 524898
rect 432438 525454 432678 525486
rect 432438 525218 432440 525454
rect 432676 525218 432678 525454
rect 432438 525134 432678 525218
rect 432438 524898 432440 525134
rect 432676 524898 432678 525134
rect 432438 524866 432678 524898
rect 433244 525454 433484 525486
rect 433244 525218 433246 525454
rect 433482 525218 433484 525454
rect 433244 525134 433484 525218
rect 433244 524898 433246 525134
rect 433482 524898 433484 525134
rect 433244 524866 433484 524898
rect 439790 525454 440030 525486
rect 439790 525218 439792 525454
rect 440028 525218 440030 525454
rect 439790 525134 440030 525218
rect 439790 524898 439792 525134
rect 440028 524898 440030 525134
rect 439790 524866 440030 524898
rect 457008 525454 457248 525486
rect 457008 525218 457010 525454
rect 457246 525218 457248 525454
rect 457008 525134 457248 525218
rect 457008 524898 457010 525134
rect 457246 524898 457248 525134
rect 457008 524866 457248 524898
rect 579288 525454 579888 525486
rect 579288 525218 579470 525454
rect 579706 525218 579888 525454
rect 579288 525134 579888 525218
rect 579288 524898 579470 525134
rect 579706 524898 579888 525134
rect 579288 524866 579888 524898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect 5200 507454 5800 507486
rect 5200 507218 5382 507454
rect 5618 507218 5800 507454
rect 5200 507134 5800 507218
rect 5200 506898 5382 507134
rect 5618 506898 5800 507134
rect 5200 506866 5800 506898
rect 127456 507454 127696 507486
rect 127456 507218 127458 507454
rect 127694 507218 127696 507454
rect 127456 507134 127696 507218
rect 127456 506898 127458 507134
rect 127694 506898 127696 507134
rect 127456 506866 127696 506898
rect 140654 507454 140894 507486
rect 140654 507218 140656 507454
rect 140892 507218 140894 507454
rect 140654 507134 140894 507218
rect 140654 506898 140656 507134
rect 140892 506898 140894 507134
rect 140654 506866 140894 506898
rect 141500 507454 141740 507486
rect 141500 507218 141502 507454
rect 141738 507218 141740 507454
rect 141500 507134 141740 507218
rect 141500 506898 141502 507134
rect 141738 506898 141740 507134
rect 141500 506866 141740 506898
rect 147286 507454 147526 507486
rect 147286 507218 147288 507454
rect 147524 507218 147526 507454
rect 147286 507134 147526 507218
rect 147286 506898 147288 507134
rect 147524 506898 147526 507134
rect 147286 506866 147526 506898
rect 149658 507454 149898 507486
rect 149658 507218 149660 507454
rect 149896 507218 149898 507454
rect 149658 507134 149898 507218
rect 149658 506898 149660 507134
rect 149896 506898 149898 507134
rect 149658 506866 149898 506898
rect 150504 507454 150744 507486
rect 150504 507218 150506 507454
rect 150742 507218 150744 507454
rect 150504 507134 150744 507218
rect 150504 506898 150506 507134
rect 150742 506898 150744 507134
rect 150504 506866 150744 506898
rect 159504 507454 159744 507486
rect 159504 507218 159506 507454
rect 159742 507218 159744 507454
rect 159504 507134 159744 507218
rect 159504 506898 159506 507134
rect 159742 506898 159744 507134
rect 159504 506866 159744 506898
rect 168504 507454 168744 507486
rect 168504 507218 168506 507454
rect 168742 507218 168744 507454
rect 168504 507134 168744 507218
rect 168504 506898 168506 507134
rect 168742 506898 168744 507134
rect 168504 506866 168744 506898
rect 177504 507454 177744 507486
rect 177504 507218 177506 507454
rect 177742 507218 177744 507454
rect 177504 507134 177744 507218
rect 177504 506898 177506 507134
rect 177742 506898 177744 507134
rect 177504 506866 177744 506898
rect 186504 507454 186744 507486
rect 186504 507218 186506 507454
rect 186742 507218 186744 507454
rect 186504 507134 186744 507218
rect 186504 506898 186506 507134
rect 186742 506898 186744 507134
rect 186504 506866 186744 506898
rect 188306 507454 188546 507486
rect 188306 507218 188308 507454
rect 188544 507218 188546 507454
rect 188306 507134 188546 507218
rect 188306 506898 188308 507134
rect 188544 506898 188546 507134
rect 188306 506866 188546 506898
rect 190678 507454 190918 507486
rect 190678 507218 190680 507454
rect 190916 507218 190918 507454
rect 190678 507134 190918 507218
rect 190678 506898 190680 507134
rect 190916 506898 190918 507134
rect 190678 506866 190918 506898
rect 191524 507454 191764 507486
rect 191524 507218 191526 507454
rect 191762 507218 191764 507454
rect 191524 507134 191764 507218
rect 191524 506898 191526 507134
rect 191762 506898 191764 507134
rect 191524 506866 191764 506898
rect 200524 507454 200764 507486
rect 200524 507218 200526 507454
rect 200762 507218 200764 507454
rect 200524 507134 200764 507218
rect 200524 506898 200526 507134
rect 200762 506898 200764 507134
rect 200524 506866 200764 506898
rect 209524 507454 209764 507486
rect 209524 507218 209526 507454
rect 209762 507218 209764 507454
rect 209524 507134 209764 507218
rect 209524 506898 209526 507134
rect 209762 506898 209764 507134
rect 209524 506866 209764 506898
rect 218524 507454 218764 507486
rect 218524 507218 218526 507454
rect 218762 507218 218764 507454
rect 218524 507134 218764 507218
rect 218524 506898 218526 507134
rect 218762 506898 218764 507134
rect 218524 506866 218764 506898
rect 227524 507454 227764 507486
rect 227524 507218 227526 507454
rect 227762 507218 227764 507454
rect 227524 507134 227764 507218
rect 227524 506898 227526 507134
rect 227762 506898 227764 507134
rect 227524 506866 227764 506898
rect 229326 507454 229566 507486
rect 229326 507218 229328 507454
rect 229564 507218 229566 507454
rect 229326 507134 229566 507218
rect 229326 506898 229328 507134
rect 229564 506898 229566 507134
rect 229326 506866 229566 506898
rect 230698 507454 230938 507486
rect 230698 507218 230700 507454
rect 230936 507218 230938 507454
rect 230698 507134 230938 507218
rect 230698 506898 230700 507134
rect 230936 506898 230938 507134
rect 230698 506866 230938 506898
rect 231544 507454 231784 507486
rect 231544 507218 231546 507454
rect 231782 507218 231784 507454
rect 231544 507134 231784 507218
rect 231544 506898 231546 507134
rect 231782 506898 231784 507134
rect 231544 506866 231784 506898
rect 240544 507454 240784 507486
rect 240544 507218 240546 507454
rect 240782 507218 240784 507454
rect 240544 507134 240784 507218
rect 240544 506898 240546 507134
rect 240782 506898 240784 507134
rect 240544 506866 240784 506898
rect 249544 507454 249784 507486
rect 249544 507218 249546 507454
rect 249782 507218 249784 507454
rect 249544 507134 249784 507218
rect 249544 506898 249546 507134
rect 249782 506898 249784 507134
rect 249544 506866 249784 506898
rect 258544 507454 258784 507486
rect 258544 507218 258546 507454
rect 258782 507218 258784 507454
rect 258544 507134 258784 507218
rect 258544 506898 258546 507134
rect 258782 506898 258784 507134
rect 258544 506866 258784 506898
rect 267544 507454 267784 507486
rect 267544 507218 267546 507454
rect 267782 507218 267784 507454
rect 267544 507134 267784 507218
rect 267544 506898 267546 507134
rect 267782 506898 267784 507134
rect 267544 506866 267784 506898
rect 269346 507454 269586 507486
rect 269346 507218 269348 507454
rect 269584 507218 269586 507454
rect 269346 507134 269586 507218
rect 269346 506898 269348 507134
rect 269584 506898 269586 507134
rect 269346 506866 269586 506898
rect 270718 507454 270958 507486
rect 270718 507218 270720 507454
rect 270956 507218 270958 507454
rect 270718 507134 270958 507218
rect 270718 506898 270720 507134
rect 270956 506898 270958 507134
rect 270718 506866 270958 506898
rect 271564 507454 271804 507486
rect 271564 507218 271566 507454
rect 271802 507218 271804 507454
rect 271564 507134 271804 507218
rect 271564 506898 271566 507134
rect 271802 506898 271804 507134
rect 271564 506866 271804 506898
rect 280564 507454 280804 507486
rect 280564 507218 280566 507454
rect 280802 507218 280804 507454
rect 280564 507134 280804 507218
rect 280564 506898 280566 507134
rect 280802 506898 280804 507134
rect 280564 506866 280804 506898
rect 289564 507454 289804 507486
rect 289564 507218 289566 507454
rect 289802 507218 289804 507454
rect 289564 507134 289804 507218
rect 289564 506898 289566 507134
rect 289802 506898 289804 507134
rect 289564 506866 289804 506898
rect 298564 507454 298804 507486
rect 298564 507218 298566 507454
rect 298802 507218 298804 507454
rect 298564 507134 298804 507218
rect 298564 506898 298566 507134
rect 298802 506898 298804 507134
rect 298564 506866 298804 506898
rect 307564 507454 307804 507486
rect 307564 507218 307566 507454
rect 307802 507218 307804 507454
rect 307564 507134 307804 507218
rect 307564 506898 307566 507134
rect 307802 506898 307804 507134
rect 307564 506866 307804 506898
rect 309366 507454 309606 507486
rect 309366 507218 309368 507454
rect 309604 507218 309606 507454
rect 309366 507134 309606 507218
rect 309366 506898 309368 507134
rect 309604 506898 309606 507134
rect 309366 506866 309606 506898
rect 311738 507454 311978 507486
rect 311738 507218 311740 507454
rect 311976 507218 311978 507454
rect 311738 507134 311978 507218
rect 311738 506898 311740 507134
rect 311976 506898 311978 507134
rect 311738 506866 311978 506898
rect 312584 507454 312824 507486
rect 312584 507218 312586 507454
rect 312822 507218 312824 507454
rect 312584 507134 312824 507218
rect 312584 506898 312586 507134
rect 312822 506898 312824 507134
rect 312584 506866 312824 506898
rect 321584 507454 321824 507486
rect 321584 507218 321586 507454
rect 321822 507218 321824 507454
rect 321584 507134 321824 507218
rect 321584 506898 321586 507134
rect 321822 506898 321824 507134
rect 321584 506866 321824 506898
rect 330584 507454 330824 507486
rect 330584 507218 330586 507454
rect 330822 507218 330824 507454
rect 330584 507134 330824 507218
rect 330584 506898 330586 507134
rect 330822 506898 330824 507134
rect 330584 506866 330824 506898
rect 339584 507454 339824 507486
rect 339584 507218 339586 507454
rect 339822 507218 339824 507454
rect 339584 507134 339824 507218
rect 339584 506898 339586 507134
rect 339822 506898 339824 507134
rect 339584 506866 339824 506898
rect 348584 507454 348824 507486
rect 348584 507218 348586 507454
rect 348822 507218 348824 507454
rect 348584 507134 348824 507218
rect 348584 506898 348586 507134
rect 348822 506898 348824 507134
rect 348584 506866 348824 506898
rect 350386 507454 350626 507486
rect 350386 507218 350388 507454
rect 350624 507218 350626 507454
rect 350386 507134 350626 507218
rect 350386 506898 350388 507134
rect 350624 506898 350626 507134
rect 350386 506866 350626 506898
rect 352758 507454 352998 507486
rect 352758 507218 352760 507454
rect 352996 507218 352998 507454
rect 352758 507134 352998 507218
rect 352758 506898 352760 507134
rect 352996 506898 352998 507134
rect 352758 506866 352998 506898
rect 353604 507454 353844 507486
rect 353604 507218 353606 507454
rect 353842 507218 353844 507454
rect 353604 507134 353844 507218
rect 353604 506898 353606 507134
rect 353842 506898 353844 507134
rect 353604 506866 353844 506898
rect 362604 507454 362844 507486
rect 362604 507218 362606 507454
rect 362842 507218 362844 507454
rect 362604 507134 362844 507218
rect 362604 506898 362606 507134
rect 362842 506898 362844 507134
rect 362604 506866 362844 506898
rect 371604 507454 371844 507486
rect 371604 507218 371606 507454
rect 371842 507218 371844 507454
rect 371604 507134 371844 507218
rect 371604 506898 371606 507134
rect 371842 506898 371844 507134
rect 371604 506866 371844 506898
rect 380604 507454 380844 507486
rect 380604 507218 380606 507454
rect 380842 507218 380844 507454
rect 380604 507134 380844 507218
rect 380604 506898 380606 507134
rect 380842 506898 380844 507134
rect 380604 506866 380844 506898
rect 389604 507454 389844 507486
rect 389604 507218 389606 507454
rect 389842 507218 389844 507454
rect 389604 507134 389844 507218
rect 389604 506898 389606 507134
rect 389842 506898 389844 507134
rect 389604 506866 389844 506898
rect 391406 507454 391646 507486
rect 391406 507218 391408 507454
rect 391644 507218 391646 507454
rect 391406 507134 391646 507218
rect 391406 506898 391408 507134
rect 391644 506898 391646 507134
rect 391406 506866 391646 506898
rect 392778 507454 393018 507486
rect 392778 507218 392780 507454
rect 393016 507218 393018 507454
rect 392778 507134 393018 507218
rect 392778 506898 392780 507134
rect 393016 506898 393018 507134
rect 392778 506866 393018 506898
rect 393624 507454 393864 507486
rect 393624 507218 393626 507454
rect 393862 507218 393864 507454
rect 393624 507134 393864 507218
rect 393624 506898 393626 507134
rect 393862 506898 393864 507134
rect 393624 506866 393864 506898
rect 402624 507454 402864 507486
rect 402624 507218 402626 507454
rect 402862 507218 402864 507454
rect 402624 507134 402864 507218
rect 402624 506898 402626 507134
rect 402862 506898 402864 507134
rect 402624 506866 402864 506898
rect 411624 507454 411864 507486
rect 411624 507218 411626 507454
rect 411862 507218 411864 507454
rect 411624 507134 411864 507218
rect 411624 506898 411626 507134
rect 411862 506898 411864 507134
rect 411624 506866 411864 506898
rect 420624 507454 420864 507486
rect 420624 507218 420626 507454
rect 420862 507218 420864 507454
rect 420624 507134 420864 507218
rect 420624 506898 420626 507134
rect 420862 506898 420864 507134
rect 420624 506866 420864 506898
rect 429624 507454 429864 507486
rect 429624 507218 429626 507454
rect 429862 507218 429864 507454
rect 429624 507134 429864 507218
rect 429624 506898 429626 507134
rect 429862 506898 429864 507134
rect 429624 506866 429864 506898
rect 431426 507454 431666 507486
rect 431426 507218 431428 507454
rect 431664 507218 431666 507454
rect 431426 507134 431666 507218
rect 431426 506898 431428 507134
rect 431664 506898 431666 507134
rect 431426 506866 431666 506898
rect 432798 507454 433038 507486
rect 432798 507218 432800 507454
rect 433036 507218 433038 507454
rect 432798 507134 433038 507218
rect 432798 506898 432800 507134
rect 433036 506898 433038 507134
rect 432798 506866 433038 506898
rect 433644 507454 433884 507486
rect 433644 507218 433646 507454
rect 433882 507218 433884 507454
rect 433644 507134 433884 507218
rect 433644 506898 433646 507134
rect 433882 506898 433884 507134
rect 433644 506866 433884 506898
rect 439430 507454 439670 507486
rect 439430 507218 439432 507454
rect 439668 507218 439670 507454
rect 439430 507134 439670 507218
rect 439430 506898 439432 507134
rect 439668 506898 439670 507134
rect 439430 506866 439670 506898
rect 456608 507454 456848 507486
rect 456608 507218 456610 507454
rect 456846 507218 456848 507454
rect 456608 507134 456848 507218
rect 456608 506898 456610 507134
rect 456846 506898 456848 507134
rect 456608 506866 456848 506898
rect 578488 507454 579088 507486
rect 578488 507218 578670 507454
rect 578906 507218 579088 507454
rect 578488 507134 579088 507218
rect 578488 506898 578670 507134
rect 578906 506898 579088 507134
rect 578488 506866 579088 506898
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 4400 489454 5000 489486
rect 4400 489218 4582 489454
rect 4818 489218 5000 489454
rect 4400 489134 5000 489218
rect 4400 488898 4582 489134
rect 4818 488898 5000 489134
rect 4400 488866 5000 488898
rect 12536 489454 12936 489486
rect 12536 489218 12618 489454
rect 12854 489218 12936 489454
rect 12536 489134 12936 489218
rect 12536 488898 12618 489134
rect 12854 488898 12936 489134
rect 12536 488866 12936 488898
rect 14040 489454 14276 489486
rect 14040 489134 14276 489218
rect 14040 488866 14276 488898
rect 23040 489454 23276 489486
rect 23040 489134 23276 489218
rect 23040 488866 23276 488898
rect 32040 489454 32276 489486
rect 32040 489134 32276 489218
rect 32040 488866 32276 488898
rect 41040 489454 41276 489486
rect 41040 489134 41276 489218
rect 41040 488866 41276 488898
rect 50040 489454 50276 489486
rect 50040 489134 50276 489218
rect 50040 488866 50276 488898
rect 59040 489454 59276 489486
rect 59040 489134 59276 489218
rect 59040 488866 59276 488898
rect 68040 489454 68276 489486
rect 68040 489134 68276 489218
rect 68040 488866 68276 488898
rect 77040 489454 77276 489486
rect 77040 489134 77276 489218
rect 77040 488866 77276 488898
rect 86040 489454 86276 489486
rect 86040 489134 86276 489218
rect 86040 488866 86276 488898
rect 95040 489454 95276 489486
rect 95040 489134 95276 489218
rect 95040 488866 95276 488898
rect 104040 489454 104276 489486
rect 104040 489134 104276 489218
rect 104040 488866 104276 488898
rect 113040 489454 113276 489486
rect 113040 489134 113276 489218
rect 113040 488866 113276 488898
rect 121144 489454 121544 489486
rect 121144 489218 121226 489454
rect 121462 489218 121544 489454
rect 121144 489134 121544 489218
rect 121144 488898 121226 489134
rect 121462 488898 121544 489134
rect 121144 488866 121544 488898
rect 127056 489454 127296 489486
rect 127056 489218 127058 489454
rect 127294 489218 127296 489454
rect 127056 489134 127296 489218
rect 127056 488898 127058 489134
rect 127294 488898 127296 489134
rect 127056 488866 127296 488898
rect 140294 489454 140534 489486
rect 140294 489218 140296 489454
rect 140532 489218 140534 489454
rect 140294 489134 140534 489218
rect 140294 488898 140296 489134
rect 140532 488898 140534 489134
rect 140294 488866 140534 488898
rect 141100 489454 141340 489486
rect 141100 489218 141102 489454
rect 141338 489218 141340 489454
rect 141100 489134 141340 489218
rect 141100 488898 141102 489134
rect 141338 488898 141340 489134
rect 141100 488866 141340 488898
rect 147646 489454 147886 489486
rect 147646 489218 147648 489454
rect 147884 489218 147886 489454
rect 147646 489134 147886 489218
rect 147646 488898 147648 489134
rect 147884 488898 147886 489134
rect 147646 488866 147886 488898
rect 149298 489454 149538 489486
rect 149298 489218 149300 489454
rect 149536 489218 149538 489454
rect 149298 489134 149538 489218
rect 149298 488898 149300 489134
rect 149536 488898 149538 489134
rect 149298 488866 149538 488898
rect 150104 489454 150344 489486
rect 150104 489218 150106 489454
rect 150342 489218 150344 489454
rect 150104 489134 150344 489218
rect 150104 488898 150106 489134
rect 150342 488898 150344 489134
rect 150104 488866 150344 488898
rect 159104 489454 159344 489486
rect 159104 489218 159106 489454
rect 159342 489218 159344 489454
rect 159104 489134 159344 489218
rect 159104 488898 159106 489134
rect 159342 488898 159344 489134
rect 159104 488866 159344 488898
rect 168104 489454 168344 489486
rect 168104 489218 168106 489454
rect 168342 489218 168344 489454
rect 168104 489134 168344 489218
rect 168104 488898 168106 489134
rect 168342 488898 168344 489134
rect 168104 488866 168344 488898
rect 177104 489454 177344 489486
rect 177104 489218 177106 489454
rect 177342 489218 177344 489454
rect 177104 489134 177344 489218
rect 177104 488898 177106 489134
rect 177342 488898 177344 489134
rect 177104 488866 177344 488898
rect 186104 489454 186344 489486
rect 186104 489218 186106 489454
rect 186342 489218 186344 489454
rect 186104 489134 186344 489218
rect 186104 488898 186106 489134
rect 186342 488898 186344 489134
rect 186104 488866 186344 488898
rect 188666 489454 188906 489486
rect 188666 489218 188668 489454
rect 188904 489218 188906 489454
rect 188666 489134 188906 489218
rect 188666 488898 188668 489134
rect 188904 488898 188906 489134
rect 188666 488866 188906 488898
rect 189766 489454 190006 489486
rect 189766 489218 189768 489454
rect 190004 489218 190006 489454
rect 189766 489134 190006 489218
rect 189766 488898 189768 489134
rect 190004 488898 190006 489134
rect 189766 488866 190006 488898
rect 190318 489454 190558 489486
rect 190318 489218 190320 489454
rect 190556 489218 190558 489454
rect 190318 489134 190558 489218
rect 190318 488898 190320 489134
rect 190556 488898 190558 489134
rect 190318 488866 190558 488898
rect 191124 489454 191364 489486
rect 191124 489218 191126 489454
rect 191362 489218 191364 489454
rect 191124 489134 191364 489218
rect 191124 488898 191126 489134
rect 191362 488898 191364 489134
rect 191124 488866 191364 488898
rect 200124 489454 200364 489486
rect 200124 489218 200126 489454
rect 200362 489218 200364 489454
rect 200124 489134 200364 489218
rect 200124 488898 200126 489134
rect 200362 488898 200364 489134
rect 200124 488866 200364 488898
rect 209124 489454 209364 489486
rect 209124 489218 209126 489454
rect 209362 489218 209364 489454
rect 209124 489134 209364 489218
rect 209124 488898 209126 489134
rect 209362 488898 209364 489134
rect 209124 488866 209364 488898
rect 218124 489454 218364 489486
rect 218124 489218 218126 489454
rect 218362 489218 218364 489454
rect 218124 489134 218364 489218
rect 218124 488898 218126 489134
rect 218362 488898 218364 489134
rect 218124 488866 218364 488898
rect 227124 489454 227364 489486
rect 227124 489218 227126 489454
rect 227362 489218 227364 489454
rect 227124 489134 227364 489218
rect 227124 488898 227126 489134
rect 227362 488898 227364 489134
rect 227124 488866 227364 488898
rect 229686 489454 229926 489486
rect 229686 489218 229688 489454
rect 229924 489218 229926 489454
rect 229686 489134 229926 489218
rect 229686 488898 229688 489134
rect 229924 488898 229926 489134
rect 229686 488866 229926 488898
rect 230338 489454 230578 489486
rect 230338 489218 230340 489454
rect 230576 489218 230578 489454
rect 230338 489134 230578 489218
rect 230338 488898 230340 489134
rect 230576 488898 230578 489134
rect 230338 488866 230578 488898
rect 231144 489454 231384 489486
rect 231144 489218 231146 489454
rect 231382 489218 231384 489454
rect 231144 489134 231384 489218
rect 231144 488898 231146 489134
rect 231382 488898 231384 489134
rect 231144 488866 231384 488898
rect 240144 489454 240384 489486
rect 240144 489218 240146 489454
rect 240382 489218 240384 489454
rect 240144 489134 240384 489218
rect 240144 488898 240146 489134
rect 240382 488898 240384 489134
rect 240144 488866 240384 488898
rect 249144 489454 249384 489486
rect 249144 489218 249146 489454
rect 249382 489218 249384 489454
rect 249144 489134 249384 489218
rect 249144 488898 249146 489134
rect 249382 488898 249384 489134
rect 249144 488866 249384 488898
rect 258144 489454 258384 489486
rect 258144 489218 258146 489454
rect 258382 489218 258384 489454
rect 258144 489134 258384 489218
rect 258144 488898 258146 489134
rect 258382 488898 258384 489134
rect 258144 488866 258384 488898
rect 267144 489454 267384 489486
rect 267144 489218 267146 489454
rect 267382 489218 267384 489454
rect 267144 489134 267384 489218
rect 267144 488898 267146 489134
rect 267382 488898 267384 489134
rect 267144 488866 267384 488898
rect 269706 489454 269946 489486
rect 269706 489218 269708 489454
rect 269944 489218 269946 489454
rect 269706 489134 269946 489218
rect 269706 488898 269708 489134
rect 269944 488898 269946 489134
rect 269706 488866 269946 488898
rect 270358 489454 270598 489486
rect 270358 489218 270360 489454
rect 270596 489218 270598 489454
rect 270358 489134 270598 489218
rect 270358 488898 270360 489134
rect 270596 488898 270598 489134
rect 270358 488866 270598 488898
rect 271164 489454 271404 489486
rect 271164 489218 271166 489454
rect 271402 489218 271404 489454
rect 271164 489134 271404 489218
rect 271164 488898 271166 489134
rect 271402 488898 271404 489134
rect 271164 488866 271404 488898
rect 280164 489454 280404 489486
rect 280164 489218 280166 489454
rect 280402 489218 280404 489454
rect 280164 489134 280404 489218
rect 280164 488898 280166 489134
rect 280402 488898 280404 489134
rect 280164 488866 280404 488898
rect 289164 489454 289404 489486
rect 289164 489218 289166 489454
rect 289402 489218 289404 489454
rect 289164 489134 289404 489218
rect 289164 488898 289166 489134
rect 289402 488898 289404 489134
rect 289164 488866 289404 488898
rect 298164 489454 298404 489486
rect 298164 489218 298166 489454
rect 298402 489218 298404 489454
rect 298164 489134 298404 489218
rect 298164 488898 298166 489134
rect 298402 488898 298404 489134
rect 298164 488866 298404 488898
rect 307164 489454 307404 489486
rect 307164 489218 307166 489454
rect 307402 489218 307404 489454
rect 307164 489134 307404 489218
rect 307164 488898 307166 489134
rect 307402 488898 307404 489134
rect 307164 488866 307404 488898
rect 309726 489454 309966 489486
rect 309726 489218 309728 489454
rect 309964 489218 309966 489454
rect 309726 489134 309966 489218
rect 309726 488898 309728 489134
rect 309964 488898 309966 489134
rect 309726 488866 309966 488898
rect 311378 489454 311618 489486
rect 311378 489218 311380 489454
rect 311616 489218 311618 489454
rect 311378 489134 311618 489218
rect 311378 488898 311380 489134
rect 311616 488898 311618 489134
rect 311378 488866 311618 488898
rect 312184 489454 312424 489486
rect 312184 489218 312186 489454
rect 312422 489218 312424 489454
rect 312184 489134 312424 489218
rect 312184 488898 312186 489134
rect 312422 488898 312424 489134
rect 312184 488866 312424 488898
rect 321184 489454 321424 489486
rect 321184 489218 321186 489454
rect 321422 489218 321424 489454
rect 321184 489134 321424 489218
rect 321184 488898 321186 489134
rect 321422 488898 321424 489134
rect 321184 488866 321424 488898
rect 330184 489454 330424 489486
rect 330184 489218 330186 489454
rect 330422 489218 330424 489454
rect 330184 489134 330424 489218
rect 330184 488898 330186 489134
rect 330422 488898 330424 489134
rect 330184 488866 330424 488898
rect 339184 489454 339424 489486
rect 339184 489218 339186 489454
rect 339422 489218 339424 489454
rect 339184 489134 339424 489218
rect 339184 488898 339186 489134
rect 339422 488898 339424 489134
rect 339184 488866 339424 488898
rect 348184 489454 348424 489486
rect 348184 489218 348186 489454
rect 348422 489218 348424 489454
rect 348184 489134 348424 489218
rect 348184 488898 348186 489134
rect 348422 488898 348424 489134
rect 348184 488866 348424 488898
rect 350746 489454 350986 489486
rect 350746 489218 350748 489454
rect 350984 489218 350986 489454
rect 350746 489134 350986 489218
rect 350746 488898 350748 489134
rect 350984 488898 350986 489134
rect 350746 488866 350986 488898
rect 352398 489454 352638 489486
rect 352398 489218 352400 489454
rect 352636 489218 352638 489454
rect 352398 489134 352638 489218
rect 352398 488898 352400 489134
rect 352636 488898 352638 489134
rect 352398 488866 352638 488898
rect 353204 489454 353444 489486
rect 353204 489218 353206 489454
rect 353442 489218 353444 489454
rect 353204 489134 353444 489218
rect 353204 488898 353206 489134
rect 353442 488898 353444 489134
rect 353204 488866 353444 488898
rect 362204 489454 362444 489486
rect 362204 489218 362206 489454
rect 362442 489218 362444 489454
rect 362204 489134 362444 489218
rect 362204 488898 362206 489134
rect 362442 488898 362444 489134
rect 362204 488866 362444 488898
rect 371204 489454 371444 489486
rect 371204 489218 371206 489454
rect 371442 489218 371444 489454
rect 371204 489134 371444 489218
rect 371204 488898 371206 489134
rect 371442 488898 371444 489134
rect 371204 488866 371444 488898
rect 380204 489454 380444 489486
rect 380204 489218 380206 489454
rect 380442 489218 380444 489454
rect 380204 489134 380444 489218
rect 380204 488898 380206 489134
rect 380442 488898 380444 489134
rect 380204 488866 380444 488898
rect 389204 489454 389444 489486
rect 389204 489218 389206 489454
rect 389442 489218 389444 489454
rect 389204 489134 389444 489218
rect 389204 488898 389206 489134
rect 389442 488898 389444 489134
rect 389204 488866 389444 488898
rect 391766 489454 392006 489486
rect 391766 489218 391768 489454
rect 392004 489218 392006 489454
rect 391766 489134 392006 489218
rect 391766 488898 391768 489134
rect 392004 488898 392006 489134
rect 391766 488866 392006 488898
rect 392418 489454 392658 489486
rect 392418 489218 392420 489454
rect 392656 489218 392658 489454
rect 392418 489134 392658 489218
rect 392418 488898 392420 489134
rect 392656 488898 392658 489134
rect 392418 488866 392658 488898
rect 393224 489454 393464 489486
rect 393224 489218 393226 489454
rect 393462 489218 393464 489454
rect 393224 489134 393464 489218
rect 393224 488898 393226 489134
rect 393462 488898 393464 489134
rect 393224 488866 393464 488898
rect 402224 489454 402464 489486
rect 402224 489218 402226 489454
rect 402462 489218 402464 489454
rect 402224 489134 402464 489218
rect 402224 488898 402226 489134
rect 402462 488898 402464 489134
rect 402224 488866 402464 488898
rect 411224 489454 411464 489486
rect 411224 489218 411226 489454
rect 411462 489218 411464 489454
rect 411224 489134 411464 489218
rect 411224 488898 411226 489134
rect 411462 488898 411464 489134
rect 411224 488866 411464 488898
rect 420224 489454 420464 489486
rect 420224 489218 420226 489454
rect 420462 489218 420464 489454
rect 420224 489134 420464 489218
rect 420224 488898 420226 489134
rect 420462 488898 420464 489134
rect 420224 488866 420464 488898
rect 429224 489454 429464 489486
rect 429224 489218 429226 489454
rect 429462 489218 429464 489454
rect 429224 489134 429464 489218
rect 429224 488898 429226 489134
rect 429462 488898 429464 489134
rect 429224 488866 429464 488898
rect 431786 489454 432026 489486
rect 431786 489218 431788 489454
rect 432024 489218 432026 489454
rect 431786 489134 432026 489218
rect 431786 488898 431788 489134
rect 432024 488898 432026 489134
rect 431786 488866 432026 488898
rect 432438 489454 432678 489486
rect 432438 489218 432440 489454
rect 432676 489218 432678 489454
rect 432438 489134 432678 489218
rect 432438 488898 432440 489134
rect 432676 488898 432678 489134
rect 432438 488866 432678 488898
rect 433244 489454 433484 489486
rect 433244 489218 433246 489454
rect 433482 489218 433484 489454
rect 433244 489134 433484 489218
rect 433244 488898 433246 489134
rect 433482 488898 433484 489134
rect 433244 488866 433484 488898
rect 439790 489454 440030 489486
rect 439790 489218 439792 489454
rect 440028 489218 440030 489454
rect 439790 489134 440030 489218
rect 439790 488898 439792 489134
rect 440028 488898 440030 489134
rect 439790 488866 440030 488898
rect 457008 489454 457248 489486
rect 457008 489218 457010 489454
rect 457246 489218 457248 489454
rect 457008 489134 457248 489218
rect 457008 488898 457010 489134
rect 457246 488898 457248 489134
rect 457008 488866 457248 488898
rect 462760 489454 463160 489486
rect 462760 489218 462842 489454
rect 463078 489218 463160 489454
rect 462760 489134 463160 489218
rect 462760 488898 462842 489134
rect 463078 488898 463160 489134
rect 462760 488866 463160 488898
rect 471028 489454 471264 489486
rect 471028 489134 471264 489218
rect 471028 488866 471264 488898
rect 480028 489454 480264 489486
rect 480028 489134 480264 489218
rect 480028 488866 480264 488898
rect 489028 489454 489264 489486
rect 489028 489134 489264 489218
rect 489028 488866 489264 488898
rect 498028 489454 498264 489486
rect 498028 489134 498264 489218
rect 498028 488866 498264 488898
rect 507028 489454 507264 489486
rect 507028 489134 507264 489218
rect 507028 488866 507264 488898
rect 516028 489454 516264 489486
rect 516028 489134 516264 489218
rect 516028 488866 516264 488898
rect 525028 489454 525264 489486
rect 525028 489134 525264 489218
rect 525028 488866 525264 488898
rect 534028 489454 534264 489486
rect 534028 489134 534264 489218
rect 534028 488866 534264 488898
rect 543028 489454 543264 489486
rect 543028 489134 543264 489218
rect 543028 488866 543264 488898
rect 552028 489454 552264 489486
rect 552028 489134 552264 489218
rect 552028 488866 552264 488898
rect 561028 489454 561264 489486
rect 561028 489134 561264 489218
rect 561028 488866 561264 488898
rect 570028 489454 570264 489486
rect 570028 489134 570264 489218
rect 570028 488866 570264 488898
rect 571368 489454 571768 489486
rect 571368 489218 571450 489454
rect 571686 489218 571768 489454
rect 571368 489134 571768 489218
rect 571368 488898 571450 489134
rect 571686 488898 571768 489134
rect 571368 488866 571768 488898
rect 579288 489454 579888 489486
rect 579288 489218 579470 489454
rect 579706 489218 579888 489454
rect 579288 489134 579888 489218
rect 579288 488898 579470 489134
rect 579706 488898 579888 489134
rect 579288 488866 579888 488898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect 5200 471454 5800 471486
rect 5200 471218 5382 471454
rect 5618 471218 5800 471454
rect 5200 471134 5800 471218
rect 5200 470898 5382 471134
rect 5618 470898 5800 471134
rect 5200 470866 5800 470898
rect 13136 471454 13536 471486
rect 13136 471218 13218 471454
rect 13454 471218 13536 471454
rect 13136 471134 13536 471218
rect 13136 470898 13218 471134
rect 13454 470898 13536 471134
rect 13136 470866 13536 470898
rect 14420 471454 14656 471486
rect 14420 471134 14656 471218
rect 14420 470866 14656 470898
rect 23420 471454 23656 471486
rect 23420 471134 23656 471218
rect 23420 470866 23656 470898
rect 32420 471454 32656 471486
rect 32420 471134 32656 471218
rect 32420 470866 32656 470898
rect 41420 471454 41656 471486
rect 41420 471134 41656 471218
rect 41420 470866 41656 470898
rect 50420 471454 50656 471486
rect 50420 471134 50656 471218
rect 50420 470866 50656 470898
rect 59420 471454 59656 471486
rect 59420 471134 59656 471218
rect 59420 470866 59656 470898
rect 68420 471454 68656 471486
rect 68420 471134 68656 471218
rect 68420 470866 68656 470898
rect 77420 471454 77656 471486
rect 77420 471134 77656 471218
rect 77420 470866 77656 470898
rect 86420 471454 86656 471486
rect 86420 471134 86656 471218
rect 86420 470866 86656 470898
rect 95420 471454 95656 471486
rect 95420 471134 95656 471218
rect 95420 470866 95656 470898
rect 104420 471454 104656 471486
rect 104420 471134 104656 471218
rect 104420 470866 104656 470898
rect 113420 471454 113656 471486
rect 113420 471134 113656 471218
rect 113420 470866 113656 470898
rect 120544 471454 120944 471486
rect 120544 471218 120626 471454
rect 120862 471218 120944 471454
rect 120544 471134 120944 471218
rect 120544 470898 120626 471134
rect 120862 470898 120944 471134
rect 120544 470866 120944 470898
rect 127456 471454 127696 471486
rect 127456 471218 127458 471454
rect 127694 471218 127696 471454
rect 127456 471134 127696 471218
rect 127456 470898 127458 471134
rect 127694 470898 127696 471134
rect 127456 470866 127696 470898
rect 140654 471454 140894 471486
rect 140654 471218 140656 471454
rect 140892 471218 140894 471454
rect 140654 471134 140894 471218
rect 140654 470898 140656 471134
rect 140892 470898 140894 471134
rect 140654 470866 140894 470898
rect 141500 471454 141740 471486
rect 141500 471218 141502 471454
rect 141738 471218 141740 471454
rect 141500 471134 141740 471218
rect 141500 470898 141502 471134
rect 141738 470898 141740 471134
rect 141500 470866 141740 470898
rect 147286 471454 147526 471486
rect 147286 471218 147288 471454
rect 147524 471218 147526 471454
rect 147286 471134 147526 471218
rect 147286 470898 147288 471134
rect 147524 470898 147526 471134
rect 147286 470866 147526 470898
rect 149658 471454 149898 471486
rect 149658 471218 149660 471454
rect 149896 471218 149898 471454
rect 149658 471134 149898 471218
rect 149658 470898 149660 471134
rect 149896 470898 149898 471134
rect 149658 470866 149898 470898
rect 150504 471454 150744 471486
rect 150504 471218 150506 471454
rect 150742 471218 150744 471454
rect 150504 471134 150744 471218
rect 150504 470898 150506 471134
rect 150742 470898 150744 471134
rect 150504 470866 150744 470898
rect 159504 471454 159744 471486
rect 159504 471218 159506 471454
rect 159742 471218 159744 471454
rect 159504 471134 159744 471218
rect 159504 470898 159506 471134
rect 159742 470898 159744 471134
rect 159504 470866 159744 470898
rect 168504 471454 168744 471486
rect 168504 471218 168506 471454
rect 168742 471218 168744 471454
rect 168504 471134 168744 471218
rect 168504 470898 168506 471134
rect 168742 470898 168744 471134
rect 168504 470866 168744 470898
rect 177504 471454 177744 471486
rect 177504 471218 177506 471454
rect 177742 471218 177744 471454
rect 177504 471134 177744 471218
rect 177504 470898 177506 471134
rect 177742 470898 177744 471134
rect 177504 470866 177744 470898
rect 186504 471454 186744 471486
rect 186504 471218 186506 471454
rect 186742 471218 186744 471454
rect 186504 471134 186744 471218
rect 186504 470898 186506 471134
rect 186742 470898 186744 471134
rect 186504 470866 186744 470898
rect 188306 471454 188546 471486
rect 188306 471218 188308 471454
rect 188544 471218 188546 471454
rect 188306 471134 188546 471218
rect 188306 470898 188308 471134
rect 188544 470898 188546 471134
rect 188306 470866 188546 470898
rect 190678 471454 190918 471486
rect 190678 471218 190680 471454
rect 190916 471218 190918 471454
rect 190678 471134 190918 471218
rect 190678 470898 190680 471134
rect 190916 470898 190918 471134
rect 190678 470866 190918 470898
rect 191524 471454 191764 471486
rect 191524 471218 191526 471454
rect 191762 471218 191764 471454
rect 191524 471134 191764 471218
rect 191524 470898 191526 471134
rect 191762 470898 191764 471134
rect 191524 470866 191764 470898
rect 200524 471454 200764 471486
rect 200524 471218 200526 471454
rect 200762 471218 200764 471454
rect 200524 471134 200764 471218
rect 200524 470898 200526 471134
rect 200762 470898 200764 471134
rect 200524 470866 200764 470898
rect 209524 471454 209764 471486
rect 209524 471218 209526 471454
rect 209762 471218 209764 471454
rect 209524 471134 209764 471218
rect 209524 470898 209526 471134
rect 209762 470898 209764 471134
rect 209524 470866 209764 470898
rect 218524 471454 218764 471486
rect 218524 471218 218526 471454
rect 218762 471218 218764 471454
rect 218524 471134 218764 471218
rect 218524 470898 218526 471134
rect 218762 470898 218764 471134
rect 218524 470866 218764 470898
rect 227524 471454 227764 471486
rect 227524 471218 227526 471454
rect 227762 471218 227764 471454
rect 227524 471134 227764 471218
rect 227524 470898 227526 471134
rect 227762 470898 227764 471134
rect 227524 470866 227764 470898
rect 229326 471454 229566 471486
rect 229326 471218 229328 471454
rect 229564 471218 229566 471454
rect 229326 471134 229566 471218
rect 229326 470898 229328 471134
rect 229564 470898 229566 471134
rect 229326 470866 229566 470898
rect 230698 471454 230938 471486
rect 230698 471218 230700 471454
rect 230936 471218 230938 471454
rect 230698 471134 230938 471218
rect 230698 470898 230700 471134
rect 230936 470898 230938 471134
rect 230698 470866 230938 470898
rect 231544 471454 231784 471486
rect 231544 471218 231546 471454
rect 231782 471218 231784 471454
rect 231544 471134 231784 471218
rect 231544 470898 231546 471134
rect 231782 470898 231784 471134
rect 231544 470866 231784 470898
rect 240544 471454 240784 471486
rect 240544 471218 240546 471454
rect 240782 471218 240784 471454
rect 240544 471134 240784 471218
rect 240544 470898 240546 471134
rect 240782 470898 240784 471134
rect 240544 470866 240784 470898
rect 249544 471454 249784 471486
rect 249544 471218 249546 471454
rect 249782 471218 249784 471454
rect 249544 471134 249784 471218
rect 249544 470898 249546 471134
rect 249782 470898 249784 471134
rect 249544 470866 249784 470898
rect 258544 471454 258784 471486
rect 258544 471218 258546 471454
rect 258782 471218 258784 471454
rect 258544 471134 258784 471218
rect 258544 470898 258546 471134
rect 258782 470898 258784 471134
rect 258544 470866 258784 470898
rect 267544 471454 267784 471486
rect 267544 471218 267546 471454
rect 267782 471218 267784 471454
rect 267544 471134 267784 471218
rect 267544 470898 267546 471134
rect 267782 470898 267784 471134
rect 267544 470866 267784 470898
rect 269346 471454 269586 471486
rect 269346 471218 269348 471454
rect 269584 471218 269586 471454
rect 269346 471134 269586 471218
rect 269346 470898 269348 471134
rect 269584 470898 269586 471134
rect 269346 470866 269586 470898
rect 270718 471454 270958 471486
rect 270718 471218 270720 471454
rect 270956 471218 270958 471454
rect 270718 471134 270958 471218
rect 270718 470898 270720 471134
rect 270956 470898 270958 471134
rect 270718 470866 270958 470898
rect 271564 471454 271804 471486
rect 271564 471218 271566 471454
rect 271802 471218 271804 471454
rect 271564 471134 271804 471218
rect 271564 470898 271566 471134
rect 271802 470898 271804 471134
rect 271564 470866 271804 470898
rect 280564 471454 280804 471486
rect 280564 471218 280566 471454
rect 280802 471218 280804 471454
rect 280564 471134 280804 471218
rect 280564 470898 280566 471134
rect 280802 470898 280804 471134
rect 280564 470866 280804 470898
rect 289564 471454 289804 471486
rect 289564 471218 289566 471454
rect 289802 471218 289804 471454
rect 289564 471134 289804 471218
rect 289564 470898 289566 471134
rect 289802 470898 289804 471134
rect 289564 470866 289804 470898
rect 298564 471454 298804 471486
rect 298564 471218 298566 471454
rect 298802 471218 298804 471454
rect 298564 471134 298804 471218
rect 298564 470898 298566 471134
rect 298802 470898 298804 471134
rect 298564 470866 298804 470898
rect 307564 471454 307804 471486
rect 307564 471218 307566 471454
rect 307802 471218 307804 471454
rect 307564 471134 307804 471218
rect 307564 470898 307566 471134
rect 307802 470898 307804 471134
rect 307564 470866 307804 470898
rect 309366 471454 309606 471486
rect 309366 471218 309368 471454
rect 309604 471218 309606 471454
rect 309366 471134 309606 471218
rect 309366 470898 309368 471134
rect 309604 470898 309606 471134
rect 309366 470866 309606 470898
rect 311738 471454 311978 471486
rect 311738 471218 311740 471454
rect 311976 471218 311978 471454
rect 311738 471134 311978 471218
rect 311738 470898 311740 471134
rect 311976 470898 311978 471134
rect 311738 470866 311978 470898
rect 312584 471454 312824 471486
rect 312584 471218 312586 471454
rect 312822 471218 312824 471454
rect 312584 471134 312824 471218
rect 312584 470898 312586 471134
rect 312822 470898 312824 471134
rect 312584 470866 312824 470898
rect 321584 471454 321824 471486
rect 321584 471218 321586 471454
rect 321822 471218 321824 471454
rect 321584 471134 321824 471218
rect 321584 470898 321586 471134
rect 321822 470898 321824 471134
rect 321584 470866 321824 470898
rect 330584 471454 330824 471486
rect 330584 471218 330586 471454
rect 330822 471218 330824 471454
rect 330584 471134 330824 471218
rect 330584 470898 330586 471134
rect 330822 470898 330824 471134
rect 330584 470866 330824 470898
rect 339584 471454 339824 471486
rect 339584 471218 339586 471454
rect 339822 471218 339824 471454
rect 339584 471134 339824 471218
rect 339584 470898 339586 471134
rect 339822 470898 339824 471134
rect 339584 470866 339824 470898
rect 348584 471454 348824 471486
rect 348584 471218 348586 471454
rect 348822 471218 348824 471454
rect 348584 471134 348824 471218
rect 348584 470898 348586 471134
rect 348822 470898 348824 471134
rect 348584 470866 348824 470898
rect 350386 471454 350626 471486
rect 350386 471218 350388 471454
rect 350624 471218 350626 471454
rect 350386 471134 350626 471218
rect 350386 470898 350388 471134
rect 350624 470898 350626 471134
rect 350386 470866 350626 470898
rect 352758 471454 352998 471486
rect 352758 471218 352760 471454
rect 352996 471218 352998 471454
rect 352758 471134 352998 471218
rect 352758 470898 352760 471134
rect 352996 470898 352998 471134
rect 352758 470866 352998 470898
rect 353604 471454 353844 471486
rect 353604 471218 353606 471454
rect 353842 471218 353844 471454
rect 353604 471134 353844 471218
rect 353604 470898 353606 471134
rect 353842 470898 353844 471134
rect 353604 470866 353844 470898
rect 362604 471454 362844 471486
rect 362604 471218 362606 471454
rect 362842 471218 362844 471454
rect 362604 471134 362844 471218
rect 362604 470898 362606 471134
rect 362842 470898 362844 471134
rect 362604 470866 362844 470898
rect 371604 471454 371844 471486
rect 371604 471218 371606 471454
rect 371842 471218 371844 471454
rect 371604 471134 371844 471218
rect 371604 470898 371606 471134
rect 371842 470898 371844 471134
rect 371604 470866 371844 470898
rect 380604 471454 380844 471486
rect 380604 471218 380606 471454
rect 380842 471218 380844 471454
rect 380604 471134 380844 471218
rect 380604 470898 380606 471134
rect 380842 470898 380844 471134
rect 380604 470866 380844 470898
rect 389604 471454 389844 471486
rect 389604 471218 389606 471454
rect 389842 471218 389844 471454
rect 389604 471134 389844 471218
rect 389604 470898 389606 471134
rect 389842 470898 389844 471134
rect 389604 470866 389844 470898
rect 391406 471454 391646 471486
rect 391406 471218 391408 471454
rect 391644 471218 391646 471454
rect 391406 471134 391646 471218
rect 391406 470898 391408 471134
rect 391644 470898 391646 471134
rect 391406 470866 391646 470898
rect 392778 471454 393018 471486
rect 392778 471218 392780 471454
rect 393016 471218 393018 471454
rect 392778 471134 393018 471218
rect 392778 470898 392780 471134
rect 393016 470898 393018 471134
rect 392778 470866 393018 470898
rect 393624 471454 393864 471486
rect 393624 471218 393626 471454
rect 393862 471218 393864 471454
rect 393624 471134 393864 471218
rect 393624 470898 393626 471134
rect 393862 470898 393864 471134
rect 393624 470866 393864 470898
rect 402624 471454 402864 471486
rect 402624 471218 402626 471454
rect 402862 471218 402864 471454
rect 402624 471134 402864 471218
rect 402624 470898 402626 471134
rect 402862 470898 402864 471134
rect 402624 470866 402864 470898
rect 411624 471454 411864 471486
rect 411624 471218 411626 471454
rect 411862 471218 411864 471454
rect 411624 471134 411864 471218
rect 411624 470898 411626 471134
rect 411862 470898 411864 471134
rect 411624 470866 411864 470898
rect 420624 471454 420864 471486
rect 420624 471218 420626 471454
rect 420862 471218 420864 471454
rect 420624 471134 420864 471218
rect 420624 470898 420626 471134
rect 420862 470898 420864 471134
rect 420624 470866 420864 470898
rect 429624 471454 429864 471486
rect 429624 471218 429626 471454
rect 429862 471218 429864 471454
rect 429624 471134 429864 471218
rect 429624 470898 429626 471134
rect 429862 470898 429864 471134
rect 429624 470866 429864 470898
rect 431426 471454 431666 471486
rect 431426 471218 431428 471454
rect 431664 471218 431666 471454
rect 431426 471134 431666 471218
rect 431426 470898 431428 471134
rect 431664 470898 431666 471134
rect 431426 470866 431666 470898
rect 432798 471454 433038 471486
rect 432798 471218 432800 471454
rect 433036 471218 433038 471454
rect 432798 471134 433038 471218
rect 432798 470898 432800 471134
rect 433036 470898 433038 471134
rect 432798 470866 433038 470898
rect 433644 471454 433884 471486
rect 433644 471218 433646 471454
rect 433882 471218 433884 471454
rect 433644 471134 433884 471218
rect 433644 470898 433646 471134
rect 433882 470898 433884 471134
rect 433644 470866 433884 470898
rect 439430 471454 439670 471486
rect 439430 471218 439432 471454
rect 439668 471218 439670 471454
rect 439430 471134 439670 471218
rect 439430 470898 439432 471134
rect 439668 470898 439670 471134
rect 439430 470866 439670 470898
rect 456608 471454 456848 471486
rect 456608 471218 456610 471454
rect 456846 471218 456848 471454
rect 456608 471134 456848 471218
rect 456608 470898 456610 471134
rect 456846 470898 456848 471134
rect 456608 470866 456848 470898
rect 463360 471454 463760 471486
rect 463360 471218 463442 471454
rect 463678 471218 463760 471454
rect 463360 471134 463760 471218
rect 463360 470898 463442 471134
rect 463678 470898 463760 471134
rect 463360 470866 463760 470898
rect 470648 471454 470884 471486
rect 470648 471134 470884 471218
rect 470648 470866 470884 470898
rect 479648 471454 479884 471486
rect 479648 471134 479884 471218
rect 479648 470866 479884 470898
rect 488648 471454 488884 471486
rect 488648 471134 488884 471218
rect 488648 470866 488884 470898
rect 497648 471454 497884 471486
rect 497648 471134 497884 471218
rect 497648 470866 497884 470898
rect 506648 471454 506884 471486
rect 506648 471134 506884 471218
rect 506648 470866 506884 470898
rect 515648 471454 515884 471486
rect 515648 471134 515884 471218
rect 515648 470866 515884 470898
rect 524648 471454 524884 471486
rect 524648 471134 524884 471218
rect 524648 470866 524884 470898
rect 533648 471454 533884 471486
rect 533648 471134 533884 471218
rect 533648 470866 533884 470898
rect 542648 471454 542884 471486
rect 542648 471134 542884 471218
rect 542648 470866 542884 470898
rect 551648 471454 551884 471486
rect 551648 471134 551884 471218
rect 551648 470866 551884 470898
rect 560648 471454 560884 471486
rect 560648 471134 560884 471218
rect 560648 470866 560884 470898
rect 569648 471454 569884 471486
rect 569648 471134 569884 471218
rect 569648 470866 569884 470898
rect 570768 471454 571168 471486
rect 570768 471218 570850 471454
rect 571086 471218 571168 471454
rect 570768 471134 571168 471218
rect 570768 470898 570850 471134
rect 571086 470898 571168 471134
rect 570768 470866 571168 470898
rect 578488 471454 579088 471486
rect 578488 471218 578670 471454
rect 578906 471218 579088 471454
rect 578488 471134 579088 471218
rect 578488 470898 578670 471134
rect 578906 470898 579088 471134
rect 578488 470866 579088 470898
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 4400 453454 5000 453486
rect 4400 453218 4582 453454
rect 4818 453218 5000 453454
rect 4400 453134 5000 453218
rect 4400 452898 4582 453134
rect 4818 452898 5000 453134
rect 4400 452866 5000 452898
rect 12536 453454 12936 453486
rect 12536 453218 12618 453454
rect 12854 453218 12936 453454
rect 12536 453134 12936 453218
rect 12536 452898 12618 453134
rect 12854 452898 12936 453134
rect 12536 452866 12936 452898
rect 14040 453454 14276 453486
rect 14040 453134 14276 453218
rect 14040 452866 14276 452898
rect 23040 453454 23276 453486
rect 23040 453134 23276 453218
rect 23040 452866 23276 452898
rect 32040 453454 32276 453486
rect 32040 453134 32276 453218
rect 32040 452866 32276 452898
rect 41040 453454 41276 453486
rect 41040 453134 41276 453218
rect 41040 452866 41276 452898
rect 50040 453454 50276 453486
rect 50040 453134 50276 453218
rect 50040 452866 50276 452898
rect 59040 453454 59276 453486
rect 59040 453134 59276 453218
rect 59040 452866 59276 452898
rect 68040 453454 68276 453486
rect 68040 453134 68276 453218
rect 68040 452866 68276 452898
rect 77040 453454 77276 453486
rect 77040 453134 77276 453218
rect 77040 452866 77276 452898
rect 86040 453454 86276 453486
rect 86040 453134 86276 453218
rect 86040 452866 86276 452898
rect 95040 453454 95276 453486
rect 95040 453134 95276 453218
rect 95040 452866 95276 452898
rect 104040 453454 104276 453486
rect 104040 453134 104276 453218
rect 104040 452866 104276 452898
rect 113040 453454 113276 453486
rect 113040 453134 113276 453218
rect 113040 452866 113276 452898
rect 121144 453454 121544 453486
rect 121144 453218 121226 453454
rect 121462 453218 121544 453454
rect 121144 453134 121544 453218
rect 121144 452898 121226 453134
rect 121462 452898 121544 453134
rect 121144 452866 121544 452898
rect 127056 453454 127296 453486
rect 127056 453218 127058 453454
rect 127294 453218 127296 453454
rect 127056 453134 127296 453218
rect 127056 452898 127058 453134
rect 127294 452898 127296 453134
rect 127056 452866 127296 452898
rect 140294 453454 140534 453486
rect 140294 453218 140296 453454
rect 140532 453218 140534 453454
rect 140294 453134 140534 453218
rect 140294 452898 140296 453134
rect 140532 452898 140534 453134
rect 140294 452866 140534 452898
rect 141100 453454 141340 453486
rect 141100 453218 141102 453454
rect 141338 453218 141340 453454
rect 141100 453134 141340 453218
rect 141100 452898 141102 453134
rect 141338 452898 141340 453134
rect 141100 452866 141340 452898
rect 147646 453454 147886 453486
rect 147646 453218 147648 453454
rect 147884 453218 147886 453454
rect 147646 453134 147886 453218
rect 147646 452898 147648 453134
rect 147884 452898 147886 453134
rect 147646 452866 147886 452898
rect 149298 453454 149538 453486
rect 149298 453218 149300 453454
rect 149536 453218 149538 453454
rect 149298 453134 149538 453218
rect 149298 452898 149300 453134
rect 149536 452898 149538 453134
rect 149298 452866 149538 452898
rect 150104 453454 150344 453486
rect 150104 453218 150106 453454
rect 150342 453218 150344 453454
rect 150104 453134 150344 453218
rect 150104 452898 150106 453134
rect 150342 452898 150344 453134
rect 150104 452866 150344 452898
rect 159104 453454 159344 453486
rect 159104 453218 159106 453454
rect 159342 453218 159344 453454
rect 159104 453134 159344 453218
rect 159104 452898 159106 453134
rect 159342 452898 159344 453134
rect 159104 452866 159344 452898
rect 168104 453454 168344 453486
rect 168104 453218 168106 453454
rect 168342 453218 168344 453454
rect 168104 453134 168344 453218
rect 168104 452898 168106 453134
rect 168342 452898 168344 453134
rect 168104 452866 168344 452898
rect 177104 453454 177344 453486
rect 177104 453218 177106 453454
rect 177342 453218 177344 453454
rect 177104 453134 177344 453218
rect 177104 452898 177106 453134
rect 177342 452898 177344 453134
rect 177104 452866 177344 452898
rect 186104 453454 186344 453486
rect 186104 453218 186106 453454
rect 186342 453218 186344 453454
rect 186104 453134 186344 453218
rect 186104 452898 186106 453134
rect 186342 452898 186344 453134
rect 186104 452866 186344 452898
rect 188666 453454 188906 453486
rect 188666 453218 188668 453454
rect 188904 453218 188906 453454
rect 188666 453134 188906 453218
rect 188666 452898 188668 453134
rect 188904 452898 188906 453134
rect 188666 452866 188906 452898
rect 190318 453454 190558 453486
rect 190318 453218 190320 453454
rect 190556 453218 190558 453454
rect 190318 453134 190558 453218
rect 190318 452898 190320 453134
rect 190556 452898 190558 453134
rect 190318 452866 190558 452898
rect 191124 453454 191364 453486
rect 191124 453218 191126 453454
rect 191362 453218 191364 453454
rect 191124 453134 191364 453218
rect 191124 452898 191126 453134
rect 191362 452898 191364 453134
rect 191124 452866 191364 452898
rect 200124 453454 200364 453486
rect 200124 453218 200126 453454
rect 200362 453218 200364 453454
rect 200124 453134 200364 453218
rect 200124 452898 200126 453134
rect 200362 452898 200364 453134
rect 200124 452866 200364 452898
rect 209124 453454 209364 453486
rect 209124 453218 209126 453454
rect 209362 453218 209364 453454
rect 209124 453134 209364 453218
rect 209124 452898 209126 453134
rect 209362 452898 209364 453134
rect 209124 452866 209364 452898
rect 218124 453454 218364 453486
rect 218124 453218 218126 453454
rect 218362 453218 218364 453454
rect 218124 453134 218364 453218
rect 218124 452898 218126 453134
rect 218362 452898 218364 453134
rect 218124 452866 218364 452898
rect 227124 453454 227364 453486
rect 227124 453218 227126 453454
rect 227362 453218 227364 453454
rect 227124 453134 227364 453218
rect 227124 452898 227126 453134
rect 227362 452898 227364 453134
rect 227124 452866 227364 452898
rect 229686 453454 229926 453486
rect 229686 453218 229688 453454
rect 229924 453218 229926 453454
rect 229686 453134 229926 453218
rect 229686 452898 229688 453134
rect 229924 452898 229926 453134
rect 229686 452866 229926 452898
rect 230338 453454 230578 453486
rect 230338 453218 230340 453454
rect 230576 453218 230578 453454
rect 230338 453134 230578 453218
rect 230338 452898 230340 453134
rect 230576 452898 230578 453134
rect 230338 452866 230578 452898
rect 231144 453454 231384 453486
rect 231144 453218 231146 453454
rect 231382 453218 231384 453454
rect 231144 453134 231384 453218
rect 231144 452898 231146 453134
rect 231382 452898 231384 453134
rect 231144 452866 231384 452898
rect 240144 453454 240384 453486
rect 240144 453218 240146 453454
rect 240382 453218 240384 453454
rect 240144 453134 240384 453218
rect 240144 452898 240146 453134
rect 240382 452898 240384 453134
rect 240144 452866 240384 452898
rect 249144 453454 249384 453486
rect 249144 453218 249146 453454
rect 249382 453218 249384 453454
rect 249144 453134 249384 453218
rect 249144 452898 249146 453134
rect 249382 452898 249384 453134
rect 249144 452866 249384 452898
rect 258144 453454 258384 453486
rect 258144 453218 258146 453454
rect 258382 453218 258384 453454
rect 258144 453134 258384 453218
rect 258144 452898 258146 453134
rect 258382 452898 258384 453134
rect 258144 452866 258384 452898
rect 267144 453454 267384 453486
rect 267144 453218 267146 453454
rect 267382 453218 267384 453454
rect 267144 453134 267384 453218
rect 267144 452898 267146 453134
rect 267382 452898 267384 453134
rect 267144 452866 267384 452898
rect 269706 453454 269946 453486
rect 269706 453218 269708 453454
rect 269944 453218 269946 453454
rect 269706 453134 269946 453218
rect 269706 452898 269708 453134
rect 269944 452898 269946 453134
rect 269706 452866 269946 452898
rect 270358 453454 270598 453486
rect 270358 453218 270360 453454
rect 270596 453218 270598 453454
rect 270358 453134 270598 453218
rect 270358 452898 270360 453134
rect 270596 452898 270598 453134
rect 270358 452866 270598 452898
rect 271164 453454 271404 453486
rect 271164 453218 271166 453454
rect 271402 453218 271404 453454
rect 271164 453134 271404 453218
rect 271164 452898 271166 453134
rect 271402 452898 271404 453134
rect 271164 452866 271404 452898
rect 280164 453454 280404 453486
rect 280164 453218 280166 453454
rect 280402 453218 280404 453454
rect 280164 453134 280404 453218
rect 280164 452898 280166 453134
rect 280402 452898 280404 453134
rect 280164 452866 280404 452898
rect 289164 453454 289404 453486
rect 289164 453218 289166 453454
rect 289402 453218 289404 453454
rect 289164 453134 289404 453218
rect 289164 452898 289166 453134
rect 289402 452898 289404 453134
rect 289164 452866 289404 452898
rect 298164 453454 298404 453486
rect 298164 453218 298166 453454
rect 298402 453218 298404 453454
rect 298164 453134 298404 453218
rect 298164 452898 298166 453134
rect 298402 452898 298404 453134
rect 298164 452866 298404 452898
rect 307164 453454 307404 453486
rect 307164 453218 307166 453454
rect 307402 453218 307404 453454
rect 307164 453134 307404 453218
rect 307164 452898 307166 453134
rect 307402 452898 307404 453134
rect 307164 452866 307404 452898
rect 309726 453454 309966 453486
rect 309726 453218 309728 453454
rect 309964 453218 309966 453454
rect 309726 453134 309966 453218
rect 309726 452898 309728 453134
rect 309964 452898 309966 453134
rect 309726 452866 309966 452898
rect 311378 453454 311618 453486
rect 311378 453218 311380 453454
rect 311616 453218 311618 453454
rect 311378 453134 311618 453218
rect 311378 452898 311380 453134
rect 311616 452898 311618 453134
rect 311378 452866 311618 452898
rect 312184 453454 312424 453486
rect 312184 453218 312186 453454
rect 312422 453218 312424 453454
rect 312184 453134 312424 453218
rect 312184 452898 312186 453134
rect 312422 452898 312424 453134
rect 312184 452866 312424 452898
rect 321184 453454 321424 453486
rect 321184 453218 321186 453454
rect 321422 453218 321424 453454
rect 321184 453134 321424 453218
rect 321184 452898 321186 453134
rect 321422 452898 321424 453134
rect 321184 452866 321424 452898
rect 330184 453454 330424 453486
rect 330184 453218 330186 453454
rect 330422 453218 330424 453454
rect 330184 453134 330424 453218
rect 330184 452898 330186 453134
rect 330422 452898 330424 453134
rect 330184 452866 330424 452898
rect 339184 453454 339424 453486
rect 339184 453218 339186 453454
rect 339422 453218 339424 453454
rect 339184 453134 339424 453218
rect 339184 452898 339186 453134
rect 339422 452898 339424 453134
rect 339184 452866 339424 452898
rect 348184 453454 348424 453486
rect 348184 453218 348186 453454
rect 348422 453218 348424 453454
rect 348184 453134 348424 453218
rect 348184 452898 348186 453134
rect 348422 452898 348424 453134
rect 348184 452866 348424 452898
rect 350746 453454 350986 453486
rect 350746 453218 350748 453454
rect 350984 453218 350986 453454
rect 350746 453134 350986 453218
rect 350746 452898 350748 453134
rect 350984 452898 350986 453134
rect 350746 452866 350986 452898
rect 352398 453454 352638 453486
rect 352398 453218 352400 453454
rect 352636 453218 352638 453454
rect 352398 453134 352638 453218
rect 352398 452898 352400 453134
rect 352636 452898 352638 453134
rect 352398 452866 352638 452898
rect 353204 453454 353444 453486
rect 353204 453218 353206 453454
rect 353442 453218 353444 453454
rect 353204 453134 353444 453218
rect 353204 452898 353206 453134
rect 353442 452898 353444 453134
rect 353204 452866 353444 452898
rect 362204 453454 362444 453486
rect 362204 453218 362206 453454
rect 362442 453218 362444 453454
rect 362204 453134 362444 453218
rect 362204 452898 362206 453134
rect 362442 452898 362444 453134
rect 362204 452866 362444 452898
rect 371204 453454 371444 453486
rect 371204 453218 371206 453454
rect 371442 453218 371444 453454
rect 371204 453134 371444 453218
rect 371204 452898 371206 453134
rect 371442 452898 371444 453134
rect 371204 452866 371444 452898
rect 380204 453454 380444 453486
rect 380204 453218 380206 453454
rect 380442 453218 380444 453454
rect 380204 453134 380444 453218
rect 380204 452898 380206 453134
rect 380442 452898 380444 453134
rect 380204 452866 380444 452898
rect 389204 453454 389444 453486
rect 389204 453218 389206 453454
rect 389442 453218 389444 453454
rect 389204 453134 389444 453218
rect 389204 452898 389206 453134
rect 389442 452898 389444 453134
rect 389204 452866 389444 452898
rect 391766 453454 392006 453486
rect 391766 453218 391768 453454
rect 392004 453218 392006 453454
rect 391766 453134 392006 453218
rect 391766 452898 391768 453134
rect 392004 452898 392006 453134
rect 391766 452866 392006 452898
rect 392418 453454 392658 453486
rect 392418 453218 392420 453454
rect 392656 453218 392658 453454
rect 392418 453134 392658 453218
rect 392418 452898 392420 453134
rect 392656 452898 392658 453134
rect 392418 452866 392658 452898
rect 393224 453454 393464 453486
rect 393224 453218 393226 453454
rect 393462 453218 393464 453454
rect 393224 453134 393464 453218
rect 393224 452898 393226 453134
rect 393462 452898 393464 453134
rect 393224 452866 393464 452898
rect 402224 453454 402464 453486
rect 402224 453218 402226 453454
rect 402462 453218 402464 453454
rect 402224 453134 402464 453218
rect 402224 452898 402226 453134
rect 402462 452898 402464 453134
rect 402224 452866 402464 452898
rect 411224 453454 411464 453486
rect 411224 453218 411226 453454
rect 411462 453218 411464 453454
rect 411224 453134 411464 453218
rect 411224 452898 411226 453134
rect 411462 452898 411464 453134
rect 411224 452866 411464 452898
rect 420224 453454 420464 453486
rect 420224 453218 420226 453454
rect 420462 453218 420464 453454
rect 420224 453134 420464 453218
rect 420224 452898 420226 453134
rect 420462 452898 420464 453134
rect 420224 452866 420464 452898
rect 429224 453454 429464 453486
rect 429224 453218 429226 453454
rect 429462 453218 429464 453454
rect 429224 453134 429464 453218
rect 429224 452898 429226 453134
rect 429462 452898 429464 453134
rect 429224 452866 429464 452898
rect 431786 453454 432026 453486
rect 431786 453218 431788 453454
rect 432024 453218 432026 453454
rect 431786 453134 432026 453218
rect 431786 452898 431788 453134
rect 432024 452898 432026 453134
rect 431786 452866 432026 452898
rect 432438 453454 432678 453486
rect 432438 453218 432440 453454
rect 432676 453218 432678 453454
rect 432438 453134 432678 453218
rect 432438 452898 432440 453134
rect 432676 452898 432678 453134
rect 432438 452866 432678 452898
rect 433244 453454 433484 453486
rect 433244 453218 433246 453454
rect 433482 453218 433484 453454
rect 433244 453134 433484 453218
rect 433244 452898 433246 453134
rect 433482 452898 433484 453134
rect 433244 452866 433484 452898
rect 439790 453454 440030 453486
rect 439790 453218 439792 453454
rect 440028 453218 440030 453454
rect 439790 453134 440030 453218
rect 439790 452898 439792 453134
rect 440028 452898 440030 453134
rect 439790 452866 440030 452898
rect 457008 453454 457248 453486
rect 457008 453218 457010 453454
rect 457246 453218 457248 453454
rect 457008 453134 457248 453218
rect 457008 452898 457010 453134
rect 457246 452898 457248 453134
rect 457008 452866 457248 452898
rect 462760 453454 463160 453486
rect 462760 453218 462842 453454
rect 463078 453218 463160 453454
rect 462760 453134 463160 453218
rect 462760 452898 462842 453134
rect 463078 452898 463160 453134
rect 462760 452866 463160 452898
rect 471028 453454 471264 453486
rect 471028 453134 471264 453218
rect 471028 452866 471264 452898
rect 480028 453454 480264 453486
rect 480028 453134 480264 453218
rect 480028 452866 480264 452898
rect 489028 453454 489264 453486
rect 489028 453134 489264 453218
rect 489028 452866 489264 452898
rect 498028 453454 498264 453486
rect 498028 453134 498264 453218
rect 498028 452866 498264 452898
rect 507028 453454 507264 453486
rect 507028 453134 507264 453218
rect 507028 452866 507264 452898
rect 516028 453454 516264 453486
rect 516028 453134 516264 453218
rect 516028 452866 516264 452898
rect 525028 453454 525264 453486
rect 525028 453134 525264 453218
rect 525028 452866 525264 452898
rect 534028 453454 534264 453486
rect 534028 453134 534264 453218
rect 534028 452866 534264 452898
rect 543028 453454 543264 453486
rect 543028 453134 543264 453218
rect 543028 452866 543264 452898
rect 552028 453454 552264 453486
rect 552028 453134 552264 453218
rect 552028 452866 552264 452898
rect 561028 453454 561264 453486
rect 561028 453134 561264 453218
rect 561028 452866 561264 452898
rect 570028 453454 570264 453486
rect 570028 453134 570264 453218
rect 570028 452866 570264 452898
rect 571368 453454 571768 453486
rect 571368 453218 571450 453454
rect 571686 453218 571768 453454
rect 571368 453134 571768 453218
rect 571368 452898 571450 453134
rect 571686 452898 571768 453134
rect 571368 452866 571768 452898
rect 579288 453454 579888 453486
rect 579288 453218 579470 453454
rect 579706 453218 579888 453454
rect 579288 453134 579888 453218
rect 579288 452898 579470 453134
rect 579706 452898 579888 453134
rect 579288 452866 579888 452898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect 5200 435454 5800 435486
rect 5200 435218 5382 435454
rect 5618 435218 5800 435454
rect 5200 435134 5800 435218
rect 5200 434898 5382 435134
rect 5618 434898 5800 435134
rect 5200 434866 5800 434898
rect 13136 435454 13536 435486
rect 13136 435218 13218 435454
rect 13454 435218 13536 435454
rect 13136 435134 13536 435218
rect 13136 434898 13218 435134
rect 13454 434898 13536 435134
rect 13136 434866 13536 434898
rect 14420 435454 14656 435486
rect 14420 435134 14656 435218
rect 14420 434866 14656 434898
rect 23420 435454 23656 435486
rect 23420 435134 23656 435218
rect 23420 434866 23656 434898
rect 32420 435454 32656 435486
rect 32420 435134 32656 435218
rect 32420 434866 32656 434898
rect 41420 435454 41656 435486
rect 41420 435134 41656 435218
rect 41420 434866 41656 434898
rect 50420 435454 50656 435486
rect 50420 435134 50656 435218
rect 50420 434866 50656 434898
rect 59420 435454 59656 435486
rect 59420 435134 59656 435218
rect 59420 434866 59656 434898
rect 68420 435454 68656 435486
rect 68420 435134 68656 435218
rect 68420 434866 68656 434898
rect 77420 435454 77656 435486
rect 77420 435134 77656 435218
rect 77420 434866 77656 434898
rect 86420 435454 86656 435486
rect 86420 435134 86656 435218
rect 86420 434866 86656 434898
rect 95420 435454 95656 435486
rect 95420 435134 95656 435218
rect 95420 434866 95656 434898
rect 104420 435454 104656 435486
rect 104420 435134 104656 435218
rect 104420 434866 104656 434898
rect 113420 435454 113656 435486
rect 113420 435134 113656 435218
rect 113420 434866 113656 434898
rect 120544 435454 120944 435486
rect 120544 435218 120626 435454
rect 120862 435218 120944 435454
rect 120544 435134 120944 435218
rect 120544 434898 120626 435134
rect 120862 434898 120944 435134
rect 120544 434866 120944 434898
rect 127456 435454 127696 435486
rect 127456 435218 127458 435454
rect 127694 435218 127696 435454
rect 127456 435134 127696 435218
rect 127456 434898 127458 435134
rect 127694 434898 127696 435134
rect 127456 434866 127696 434898
rect 140654 435454 140894 435486
rect 140654 435218 140656 435454
rect 140892 435218 140894 435454
rect 140654 435134 140894 435218
rect 140654 434898 140656 435134
rect 140892 434898 140894 435134
rect 140654 434866 140894 434898
rect 147286 435454 147526 435486
rect 147286 435218 147288 435454
rect 147524 435218 147526 435454
rect 147286 435134 147526 435218
rect 147286 434898 147288 435134
rect 147524 434898 147526 435134
rect 147286 434866 147526 434898
rect 149658 435454 149898 435486
rect 149658 435218 149660 435454
rect 149896 435218 149898 435454
rect 149658 435134 149898 435218
rect 149658 434898 149660 435134
rect 149896 434898 149898 435134
rect 149658 434866 149898 434898
rect 150504 435454 150744 435486
rect 150504 435218 150506 435454
rect 150742 435218 150744 435454
rect 150504 435134 150744 435218
rect 150504 434898 150506 435134
rect 150742 434898 150744 435134
rect 150504 434866 150744 434898
rect 159504 435454 159744 435486
rect 159504 435218 159506 435454
rect 159742 435218 159744 435454
rect 159504 435134 159744 435218
rect 159504 434898 159506 435134
rect 159742 434898 159744 435134
rect 159504 434866 159744 434898
rect 168504 435454 168744 435486
rect 168504 435218 168506 435454
rect 168742 435218 168744 435454
rect 168504 435134 168744 435218
rect 168504 434898 168506 435134
rect 168742 434898 168744 435134
rect 168504 434866 168744 434898
rect 177504 435454 177744 435486
rect 177504 435218 177506 435454
rect 177742 435218 177744 435454
rect 177504 435134 177744 435218
rect 177504 434898 177506 435134
rect 177742 434898 177744 435134
rect 177504 434866 177744 434898
rect 186504 435454 186744 435486
rect 186504 435218 186506 435454
rect 186742 435218 186744 435454
rect 186504 435134 186744 435218
rect 186504 434898 186506 435134
rect 186742 434898 186744 435134
rect 186504 434866 186744 434898
rect 188306 435454 188546 435486
rect 188306 435218 188308 435454
rect 188544 435218 188546 435454
rect 188306 435134 188546 435218
rect 188306 434898 188308 435134
rect 188544 434898 188546 435134
rect 188306 434866 188546 434898
rect 190678 435454 190918 435486
rect 190678 435218 190680 435454
rect 190916 435218 190918 435454
rect 190678 435134 190918 435218
rect 190678 434898 190680 435134
rect 190916 434898 190918 435134
rect 190678 434866 190918 434898
rect 229326 435454 229566 435486
rect 229326 435218 229328 435454
rect 229564 435218 229566 435454
rect 229326 435134 229566 435218
rect 229326 434898 229328 435134
rect 229564 434898 229566 435134
rect 229326 434866 229566 434898
rect 230698 435454 230938 435486
rect 230698 435218 230700 435454
rect 230936 435218 230938 435454
rect 230698 435134 230938 435218
rect 230698 434898 230700 435134
rect 230936 434898 230938 435134
rect 230698 434866 230938 434898
rect 269346 435454 269586 435486
rect 269346 435218 269348 435454
rect 269584 435218 269586 435454
rect 269346 435134 269586 435218
rect 269346 434898 269348 435134
rect 269584 434898 269586 435134
rect 269346 434866 269586 434898
rect 270718 435454 270958 435486
rect 270718 435218 270720 435454
rect 270956 435218 270958 435454
rect 270718 435134 270958 435218
rect 270718 434898 270720 435134
rect 270956 434898 270958 435134
rect 270718 434866 270958 434898
rect 309366 435454 309606 435486
rect 309366 435218 309368 435454
rect 309604 435218 309606 435454
rect 309366 435134 309606 435218
rect 309366 434898 309368 435134
rect 309604 434898 309606 435134
rect 309366 434866 309606 434898
rect 311738 435454 311978 435486
rect 311738 435218 311740 435454
rect 311976 435218 311978 435454
rect 311738 435134 311978 435218
rect 311738 434898 311740 435134
rect 311976 434898 311978 435134
rect 311738 434866 311978 434898
rect 312584 435454 312824 435486
rect 312584 435218 312586 435454
rect 312822 435218 312824 435454
rect 312584 435134 312824 435218
rect 312584 434898 312586 435134
rect 312822 434898 312824 435134
rect 312584 434866 312824 434898
rect 321584 435454 321824 435486
rect 321584 435218 321586 435454
rect 321822 435218 321824 435454
rect 321584 435134 321824 435218
rect 321584 434898 321586 435134
rect 321822 434898 321824 435134
rect 321584 434866 321824 434898
rect 330584 435454 330824 435486
rect 330584 435218 330586 435454
rect 330822 435218 330824 435454
rect 330584 435134 330824 435218
rect 330584 434898 330586 435134
rect 330822 434898 330824 435134
rect 330584 434866 330824 434898
rect 339584 435454 339824 435486
rect 339584 435218 339586 435454
rect 339822 435218 339824 435454
rect 339584 435134 339824 435218
rect 339584 434898 339586 435134
rect 339822 434898 339824 435134
rect 339584 434866 339824 434898
rect 348584 435454 348824 435486
rect 348584 435218 348586 435454
rect 348822 435218 348824 435454
rect 348584 435134 348824 435218
rect 348584 434898 348586 435134
rect 348822 434898 348824 435134
rect 348584 434866 348824 434898
rect 350386 435454 350626 435486
rect 350386 435218 350388 435454
rect 350624 435218 350626 435454
rect 350386 435134 350626 435218
rect 350386 434898 350388 435134
rect 350624 434898 350626 435134
rect 350386 434866 350626 434898
rect 352758 435454 352998 435486
rect 352758 435218 352760 435454
rect 352996 435218 352998 435454
rect 352758 435134 352998 435218
rect 352758 434898 352760 435134
rect 352996 434898 352998 435134
rect 352758 434866 352998 434898
rect 391406 435454 391646 435486
rect 391406 435218 391408 435454
rect 391644 435218 391646 435454
rect 391406 435134 391646 435218
rect 391406 434898 391408 435134
rect 391644 434898 391646 435134
rect 391406 434866 391646 434898
rect 392778 435454 393018 435486
rect 392778 435218 392780 435454
rect 393016 435218 393018 435454
rect 392778 435134 393018 435218
rect 392778 434898 392780 435134
rect 393016 434898 393018 435134
rect 392778 434866 393018 434898
rect 431426 435454 431666 435486
rect 431426 435218 431428 435454
rect 431664 435218 431666 435454
rect 431426 435134 431666 435218
rect 431426 434898 431428 435134
rect 431664 434898 431666 435134
rect 431426 434866 431666 434898
rect 432798 435454 433038 435486
rect 432798 435218 432800 435454
rect 433036 435218 433038 435454
rect 432798 435134 433038 435218
rect 432798 434898 432800 435134
rect 433036 434898 433038 435134
rect 432798 434866 433038 434898
rect 439430 435454 439670 435486
rect 439430 435218 439432 435454
rect 439668 435218 439670 435454
rect 439430 435134 439670 435218
rect 439430 434898 439432 435134
rect 439668 434898 439670 435134
rect 439430 434866 439670 434898
rect 456608 435454 456848 435486
rect 456608 435218 456610 435454
rect 456846 435218 456848 435454
rect 456608 435134 456848 435218
rect 456608 434898 456610 435134
rect 456846 434898 456848 435134
rect 456608 434866 456848 434898
rect 463360 435454 463760 435486
rect 463360 435218 463442 435454
rect 463678 435218 463760 435454
rect 463360 435134 463760 435218
rect 463360 434898 463442 435134
rect 463678 434898 463760 435134
rect 463360 434866 463760 434898
rect 470648 435454 470884 435486
rect 470648 435134 470884 435218
rect 470648 434866 470884 434898
rect 479648 435454 479884 435486
rect 479648 435134 479884 435218
rect 479648 434866 479884 434898
rect 488648 435454 488884 435486
rect 488648 435134 488884 435218
rect 488648 434866 488884 434898
rect 497648 435454 497884 435486
rect 497648 435134 497884 435218
rect 497648 434866 497884 434898
rect 506648 435454 506884 435486
rect 506648 435134 506884 435218
rect 506648 434866 506884 434898
rect 515648 435454 515884 435486
rect 515648 435134 515884 435218
rect 515648 434866 515884 434898
rect 524648 435454 524884 435486
rect 524648 435134 524884 435218
rect 524648 434866 524884 434898
rect 533648 435454 533884 435486
rect 533648 435134 533884 435218
rect 533648 434866 533884 434898
rect 542648 435454 542884 435486
rect 542648 435134 542884 435218
rect 542648 434866 542884 434898
rect 551648 435454 551884 435486
rect 551648 435134 551884 435218
rect 551648 434866 551884 434898
rect 560648 435454 560884 435486
rect 560648 435134 560884 435218
rect 560648 434866 560884 434898
rect 569648 435454 569884 435486
rect 569648 435134 569884 435218
rect 569648 434866 569884 434898
rect 570768 435454 571168 435486
rect 570768 435218 570850 435454
rect 571086 435218 571168 435454
rect 570768 435134 571168 435218
rect 570768 434898 570850 435134
rect 571086 434898 571168 435134
rect 570768 434866 571168 434898
rect 578488 435454 579088 435486
rect 578488 435218 578670 435454
rect 578906 435218 579088 435454
rect 578488 435134 579088 435218
rect 578488 434898 578670 435134
rect 578906 434898 579088 435134
rect 578488 434866 579088 434898
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 4400 417454 5000 417486
rect 4400 417218 4582 417454
rect 4818 417218 5000 417454
rect 4400 417134 5000 417218
rect 4400 416898 4582 417134
rect 4818 416898 5000 417134
rect 4400 416866 5000 416898
rect 12536 417454 12936 417486
rect 12536 417218 12618 417454
rect 12854 417218 12936 417454
rect 12536 417134 12936 417218
rect 12536 416898 12618 417134
rect 12854 416898 12936 417134
rect 12536 416866 12936 416898
rect 14040 417454 14276 417486
rect 14040 417134 14276 417218
rect 14040 416866 14276 416898
rect 23040 417454 23276 417486
rect 23040 417134 23276 417218
rect 23040 416866 23276 416898
rect 32040 417454 32276 417486
rect 32040 417134 32276 417218
rect 32040 416866 32276 416898
rect 41040 417454 41276 417486
rect 41040 417134 41276 417218
rect 41040 416866 41276 416898
rect 50040 417454 50276 417486
rect 50040 417134 50276 417218
rect 50040 416866 50276 416898
rect 59040 417454 59276 417486
rect 59040 417134 59276 417218
rect 59040 416866 59276 416898
rect 68040 417454 68276 417486
rect 68040 417134 68276 417218
rect 68040 416866 68276 416898
rect 77040 417454 77276 417486
rect 77040 417134 77276 417218
rect 77040 416866 77276 416898
rect 86040 417454 86276 417486
rect 86040 417134 86276 417218
rect 86040 416866 86276 416898
rect 95040 417454 95276 417486
rect 95040 417134 95276 417218
rect 95040 416866 95276 416898
rect 104040 417454 104276 417486
rect 104040 417134 104276 417218
rect 104040 416866 104276 416898
rect 113040 417454 113276 417486
rect 113040 417134 113276 417218
rect 113040 416866 113276 416898
rect 121144 417454 121544 417486
rect 121144 417218 121226 417454
rect 121462 417218 121544 417454
rect 121144 417134 121544 417218
rect 121144 416898 121226 417134
rect 121462 416898 121544 417134
rect 121144 416866 121544 416898
rect 127056 417454 127296 417486
rect 127056 417218 127058 417454
rect 127294 417218 127296 417454
rect 127056 417134 127296 417218
rect 127056 416898 127058 417134
rect 127294 416898 127296 417134
rect 127056 416866 127296 416898
rect 140294 417454 140534 417486
rect 140294 417218 140296 417454
rect 140532 417218 140534 417454
rect 140294 417134 140534 417218
rect 140294 416898 140296 417134
rect 140532 416898 140534 417134
rect 140294 416866 140534 416898
rect 141100 417454 141340 417486
rect 141100 417218 141102 417454
rect 141338 417218 141340 417454
rect 141100 417134 141340 417218
rect 141100 416898 141102 417134
rect 141338 416898 141340 417134
rect 141100 416866 141340 416898
rect 147646 417454 147886 417486
rect 147646 417218 147648 417454
rect 147884 417218 147886 417454
rect 147646 417134 147886 417218
rect 147646 416898 147648 417134
rect 147884 416898 147886 417134
rect 147646 416866 147886 416898
rect 149298 417454 149538 417486
rect 149298 417218 149300 417454
rect 149536 417218 149538 417454
rect 149298 417134 149538 417218
rect 149298 416898 149300 417134
rect 149536 416898 149538 417134
rect 149298 416866 149538 416898
rect 150104 417454 150344 417486
rect 150104 417218 150106 417454
rect 150342 417218 150344 417454
rect 150104 417134 150344 417218
rect 150104 416898 150106 417134
rect 150342 416898 150344 417134
rect 150104 416866 150344 416898
rect 159104 417454 159344 417486
rect 159104 417218 159106 417454
rect 159342 417218 159344 417454
rect 159104 417134 159344 417218
rect 159104 416898 159106 417134
rect 159342 416898 159344 417134
rect 159104 416866 159344 416898
rect 168104 417454 168344 417486
rect 168104 417218 168106 417454
rect 168342 417218 168344 417454
rect 168104 417134 168344 417218
rect 168104 416898 168106 417134
rect 168342 416898 168344 417134
rect 168104 416866 168344 416898
rect 177104 417454 177344 417486
rect 177104 417218 177106 417454
rect 177342 417218 177344 417454
rect 177104 417134 177344 417218
rect 177104 416898 177106 417134
rect 177342 416898 177344 417134
rect 177104 416866 177344 416898
rect 186104 417454 186344 417486
rect 186104 417218 186106 417454
rect 186342 417218 186344 417454
rect 186104 417134 186344 417218
rect 186104 416898 186106 417134
rect 186342 416898 186344 417134
rect 186104 416866 186344 416898
rect 188666 417454 188906 417486
rect 188666 417218 188668 417454
rect 188904 417218 188906 417454
rect 188666 417134 188906 417218
rect 188666 416898 188668 417134
rect 188904 416898 188906 417134
rect 188666 416866 188906 416898
rect 189766 417454 190006 417486
rect 189766 417218 189768 417454
rect 190004 417218 190006 417454
rect 189766 417134 190006 417218
rect 189766 416898 189768 417134
rect 190004 416898 190006 417134
rect 189766 416866 190006 416898
rect 190318 417454 190558 417486
rect 190318 417218 190320 417454
rect 190556 417218 190558 417454
rect 190318 417134 190558 417218
rect 190318 416898 190320 417134
rect 190556 416898 190558 417134
rect 190318 416866 190558 416898
rect 191124 417454 191364 417486
rect 191124 417218 191126 417454
rect 191362 417218 191364 417454
rect 191124 417134 191364 417218
rect 191124 416898 191126 417134
rect 191362 416898 191364 417134
rect 191124 416866 191364 416898
rect 200124 417454 200364 417486
rect 200124 417218 200126 417454
rect 200362 417218 200364 417454
rect 200124 417134 200364 417218
rect 200124 416898 200126 417134
rect 200362 416898 200364 417134
rect 200124 416866 200364 416898
rect 209124 417454 209364 417486
rect 209124 417218 209126 417454
rect 209362 417218 209364 417454
rect 209124 417134 209364 417218
rect 209124 416898 209126 417134
rect 209362 416898 209364 417134
rect 209124 416866 209364 416898
rect 218124 417454 218364 417486
rect 218124 417218 218126 417454
rect 218362 417218 218364 417454
rect 218124 417134 218364 417218
rect 218124 416898 218126 417134
rect 218362 416898 218364 417134
rect 218124 416866 218364 416898
rect 227124 417454 227364 417486
rect 227124 417218 227126 417454
rect 227362 417218 227364 417454
rect 227124 417134 227364 417218
rect 227124 416898 227126 417134
rect 227362 416898 227364 417134
rect 227124 416866 227364 416898
rect 229686 417454 229926 417486
rect 229686 417218 229688 417454
rect 229924 417218 229926 417454
rect 229686 417134 229926 417218
rect 229686 416898 229688 417134
rect 229924 416898 229926 417134
rect 229686 416866 229926 416898
rect 230338 417454 230578 417486
rect 230338 417218 230340 417454
rect 230576 417218 230578 417454
rect 230338 417134 230578 417218
rect 230338 416898 230340 417134
rect 230576 416898 230578 417134
rect 230338 416866 230578 416898
rect 231144 417454 231384 417486
rect 231144 417218 231146 417454
rect 231382 417218 231384 417454
rect 231144 417134 231384 417218
rect 231144 416898 231146 417134
rect 231382 416898 231384 417134
rect 231144 416866 231384 416898
rect 240144 417454 240384 417486
rect 240144 417218 240146 417454
rect 240382 417218 240384 417454
rect 240144 417134 240384 417218
rect 240144 416898 240146 417134
rect 240382 416898 240384 417134
rect 240144 416866 240384 416898
rect 249144 417454 249384 417486
rect 249144 417218 249146 417454
rect 249382 417218 249384 417454
rect 249144 417134 249384 417218
rect 249144 416898 249146 417134
rect 249382 416898 249384 417134
rect 249144 416866 249384 416898
rect 258144 417454 258384 417486
rect 258144 417218 258146 417454
rect 258382 417218 258384 417454
rect 258144 417134 258384 417218
rect 258144 416898 258146 417134
rect 258382 416898 258384 417134
rect 258144 416866 258384 416898
rect 267144 417454 267384 417486
rect 267144 417218 267146 417454
rect 267382 417218 267384 417454
rect 267144 417134 267384 417218
rect 267144 416898 267146 417134
rect 267382 416898 267384 417134
rect 267144 416866 267384 416898
rect 269706 417454 269946 417486
rect 269706 417218 269708 417454
rect 269944 417218 269946 417454
rect 269706 417134 269946 417218
rect 269706 416898 269708 417134
rect 269944 416898 269946 417134
rect 269706 416866 269946 416898
rect 270358 417454 270598 417486
rect 270358 417218 270360 417454
rect 270596 417218 270598 417454
rect 270358 417134 270598 417218
rect 270358 416898 270360 417134
rect 270596 416898 270598 417134
rect 270358 416866 270598 416898
rect 271164 417454 271404 417486
rect 271164 417218 271166 417454
rect 271402 417218 271404 417454
rect 271164 417134 271404 417218
rect 271164 416898 271166 417134
rect 271402 416898 271404 417134
rect 271164 416866 271404 416898
rect 280164 417454 280404 417486
rect 280164 417218 280166 417454
rect 280402 417218 280404 417454
rect 280164 417134 280404 417218
rect 280164 416898 280166 417134
rect 280402 416898 280404 417134
rect 280164 416866 280404 416898
rect 289164 417454 289404 417486
rect 289164 417218 289166 417454
rect 289402 417218 289404 417454
rect 289164 417134 289404 417218
rect 289164 416898 289166 417134
rect 289402 416898 289404 417134
rect 289164 416866 289404 416898
rect 298164 417454 298404 417486
rect 298164 417218 298166 417454
rect 298402 417218 298404 417454
rect 298164 417134 298404 417218
rect 298164 416898 298166 417134
rect 298402 416898 298404 417134
rect 298164 416866 298404 416898
rect 307164 417454 307404 417486
rect 307164 417218 307166 417454
rect 307402 417218 307404 417454
rect 307164 417134 307404 417218
rect 307164 416898 307166 417134
rect 307402 416898 307404 417134
rect 307164 416866 307404 416898
rect 309726 417454 309966 417486
rect 309726 417218 309728 417454
rect 309964 417218 309966 417454
rect 309726 417134 309966 417218
rect 309726 416898 309728 417134
rect 309964 416898 309966 417134
rect 309726 416866 309966 416898
rect 311378 417454 311618 417486
rect 311378 417218 311380 417454
rect 311616 417218 311618 417454
rect 311378 417134 311618 417218
rect 311378 416898 311380 417134
rect 311616 416898 311618 417134
rect 311378 416866 311618 416898
rect 312184 417454 312424 417486
rect 312184 417218 312186 417454
rect 312422 417218 312424 417454
rect 312184 417134 312424 417218
rect 312184 416898 312186 417134
rect 312422 416898 312424 417134
rect 312184 416866 312424 416898
rect 321184 417454 321424 417486
rect 321184 417218 321186 417454
rect 321422 417218 321424 417454
rect 321184 417134 321424 417218
rect 321184 416898 321186 417134
rect 321422 416898 321424 417134
rect 321184 416866 321424 416898
rect 330184 417454 330424 417486
rect 330184 417218 330186 417454
rect 330422 417218 330424 417454
rect 330184 417134 330424 417218
rect 330184 416898 330186 417134
rect 330422 416898 330424 417134
rect 330184 416866 330424 416898
rect 339184 417454 339424 417486
rect 339184 417218 339186 417454
rect 339422 417218 339424 417454
rect 339184 417134 339424 417218
rect 339184 416898 339186 417134
rect 339422 416898 339424 417134
rect 339184 416866 339424 416898
rect 348184 417454 348424 417486
rect 348184 417218 348186 417454
rect 348422 417218 348424 417454
rect 348184 417134 348424 417218
rect 348184 416898 348186 417134
rect 348422 416898 348424 417134
rect 348184 416866 348424 416898
rect 350746 417454 350986 417486
rect 350746 417218 350748 417454
rect 350984 417218 350986 417454
rect 350746 417134 350986 417218
rect 350746 416898 350748 417134
rect 350984 416898 350986 417134
rect 350746 416866 350986 416898
rect 352398 417454 352638 417486
rect 352398 417218 352400 417454
rect 352636 417218 352638 417454
rect 352398 417134 352638 417218
rect 352398 416898 352400 417134
rect 352636 416898 352638 417134
rect 352398 416866 352638 416898
rect 353204 417454 353444 417486
rect 353204 417218 353206 417454
rect 353442 417218 353444 417454
rect 353204 417134 353444 417218
rect 353204 416898 353206 417134
rect 353442 416898 353444 417134
rect 353204 416866 353444 416898
rect 362204 417454 362444 417486
rect 362204 417218 362206 417454
rect 362442 417218 362444 417454
rect 362204 417134 362444 417218
rect 362204 416898 362206 417134
rect 362442 416898 362444 417134
rect 362204 416866 362444 416898
rect 371204 417454 371444 417486
rect 371204 417218 371206 417454
rect 371442 417218 371444 417454
rect 371204 417134 371444 417218
rect 371204 416898 371206 417134
rect 371442 416898 371444 417134
rect 371204 416866 371444 416898
rect 380204 417454 380444 417486
rect 380204 417218 380206 417454
rect 380442 417218 380444 417454
rect 380204 417134 380444 417218
rect 380204 416898 380206 417134
rect 380442 416898 380444 417134
rect 380204 416866 380444 416898
rect 389204 417454 389444 417486
rect 389204 417218 389206 417454
rect 389442 417218 389444 417454
rect 389204 417134 389444 417218
rect 389204 416898 389206 417134
rect 389442 416898 389444 417134
rect 389204 416866 389444 416898
rect 391766 417454 392006 417486
rect 391766 417218 391768 417454
rect 392004 417218 392006 417454
rect 391766 417134 392006 417218
rect 391766 416898 391768 417134
rect 392004 416898 392006 417134
rect 391766 416866 392006 416898
rect 392418 417454 392658 417486
rect 392418 417218 392420 417454
rect 392656 417218 392658 417454
rect 392418 417134 392658 417218
rect 392418 416898 392420 417134
rect 392656 416898 392658 417134
rect 392418 416866 392658 416898
rect 393224 417454 393464 417486
rect 393224 417218 393226 417454
rect 393462 417218 393464 417454
rect 393224 417134 393464 417218
rect 393224 416898 393226 417134
rect 393462 416898 393464 417134
rect 393224 416866 393464 416898
rect 402224 417454 402464 417486
rect 402224 417218 402226 417454
rect 402462 417218 402464 417454
rect 402224 417134 402464 417218
rect 402224 416898 402226 417134
rect 402462 416898 402464 417134
rect 402224 416866 402464 416898
rect 411224 417454 411464 417486
rect 411224 417218 411226 417454
rect 411462 417218 411464 417454
rect 411224 417134 411464 417218
rect 411224 416898 411226 417134
rect 411462 416898 411464 417134
rect 411224 416866 411464 416898
rect 420224 417454 420464 417486
rect 420224 417218 420226 417454
rect 420462 417218 420464 417454
rect 420224 417134 420464 417218
rect 420224 416898 420226 417134
rect 420462 416898 420464 417134
rect 420224 416866 420464 416898
rect 429224 417454 429464 417486
rect 429224 417218 429226 417454
rect 429462 417218 429464 417454
rect 429224 417134 429464 417218
rect 429224 416898 429226 417134
rect 429462 416898 429464 417134
rect 429224 416866 429464 416898
rect 431786 417454 432026 417486
rect 431786 417218 431788 417454
rect 432024 417218 432026 417454
rect 431786 417134 432026 417218
rect 431786 416898 431788 417134
rect 432024 416898 432026 417134
rect 431786 416866 432026 416898
rect 432438 417454 432678 417486
rect 432438 417218 432440 417454
rect 432676 417218 432678 417454
rect 432438 417134 432678 417218
rect 432438 416898 432440 417134
rect 432676 416898 432678 417134
rect 432438 416866 432678 416898
rect 433244 417454 433484 417486
rect 433244 417218 433246 417454
rect 433482 417218 433484 417454
rect 433244 417134 433484 417218
rect 433244 416898 433246 417134
rect 433482 416898 433484 417134
rect 433244 416866 433484 416898
rect 439790 417454 440030 417486
rect 439790 417218 439792 417454
rect 440028 417218 440030 417454
rect 439790 417134 440030 417218
rect 439790 416898 439792 417134
rect 440028 416898 440030 417134
rect 439790 416866 440030 416898
rect 457008 417454 457248 417486
rect 457008 417218 457010 417454
rect 457246 417218 457248 417454
rect 457008 417134 457248 417218
rect 457008 416898 457010 417134
rect 457246 416898 457248 417134
rect 457008 416866 457248 416898
rect 462760 417454 463160 417486
rect 462760 417218 462842 417454
rect 463078 417218 463160 417454
rect 462760 417134 463160 417218
rect 462760 416898 462842 417134
rect 463078 416898 463160 417134
rect 462760 416866 463160 416898
rect 471028 417454 471264 417486
rect 471028 417134 471264 417218
rect 471028 416866 471264 416898
rect 480028 417454 480264 417486
rect 480028 417134 480264 417218
rect 480028 416866 480264 416898
rect 489028 417454 489264 417486
rect 489028 417134 489264 417218
rect 489028 416866 489264 416898
rect 498028 417454 498264 417486
rect 498028 417134 498264 417218
rect 498028 416866 498264 416898
rect 507028 417454 507264 417486
rect 507028 417134 507264 417218
rect 507028 416866 507264 416898
rect 516028 417454 516264 417486
rect 516028 417134 516264 417218
rect 516028 416866 516264 416898
rect 525028 417454 525264 417486
rect 525028 417134 525264 417218
rect 525028 416866 525264 416898
rect 534028 417454 534264 417486
rect 534028 417134 534264 417218
rect 534028 416866 534264 416898
rect 543028 417454 543264 417486
rect 543028 417134 543264 417218
rect 543028 416866 543264 416898
rect 552028 417454 552264 417486
rect 552028 417134 552264 417218
rect 552028 416866 552264 416898
rect 561028 417454 561264 417486
rect 561028 417134 561264 417218
rect 561028 416866 561264 416898
rect 570028 417454 570264 417486
rect 570028 417134 570264 417218
rect 570028 416866 570264 416898
rect 571368 417454 571768 417486
rect 571368 417218 571450 417454
rect 571686 417218 571768 417454
rect 571368 417134 571768 417218
rect 571368 416898 571450 417134
rect 571686 416898 571768 417134
rect 571368 416866 571768 416898
rect 579288 417454 579888 417486
rect 579288 417218 579470 417454
rect 579706 417218 579888 417454
rect 579288 417134 579888 417218
rect 579288 416898 579470 417134
rect 579706 416898 579888 417134
rect 579288 416866 579888 416898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect 5200 399454 5800 399486
rect 5200 399218 5382 399454
rect 5618 399218 5800 399454
rect 5200 399134 5800 399218
rect 5200 398898 5382 399134
rect 5618 398898 5800 399134
rect 5200 398866 5800 398898
rect 13136 399454 13536 399486
rect 13136 399218 13218 399454
rect 13454 399218 13536 399454
rect 13136 399134 13536 399218
rect 13136 398898 13218 399134
rect 13454 398898 13536 399134
rect 13136 398866 13536 398898
rect 14420 399454 14656 399486
rect 14420 399134 14656 399218
rect 14420 398866 14656 398898
rect 23420 399454 23656 399486
rect 23420 399134 23656 399218
rect 23420 398866 23656 398898
rect 32420 399454 32656 399486
rect 32420 399134 32656 399218
rect 32420 398866 32656 398898
rect 41420 399454 41656 399486
rect 41420 399134 41656 399218
rect 41420 398866 41656 398898
rect 50420 399454 50656 399486
rect 50420 399134 50656 399218
rect 50420 398866 50656 398898
rect 59420 399454 59656 399486
rect 59420 399134 59656 399218
rect 59420 398866 59656 398898
rect 68420 399454 68656 399486
rect 68420 399134 68656 399218
rect 68420 398866 68656 398898
rect 77420 399454 77656 399486
rect 77420 399134 77656 399218
rect 77420 398866 77656 398898
rect 86420 399454 86656 399486
rect 86420 399134 86656 399218
rect 86420 398866 86656 398898
rect 95420 399454 95656 399486
rect 95420 399134 95656 399218
rect 95420 398866 95656 398898
rect 104420 399454 104656 399486
rect 104420 399134 104656 399218
rect 104420 398866 104656 398898
rect 113420 399454 113656 399486
rect 113420 399134 113656 399218
rect 113420 398866 113656 398898
rect 120544 399454 120944 399486
rect 120544 399218 120626 399454
rect 120862 399218 120944 399454
rect 120544 399134 120944 399218
rect 120544 398898 120626 399134
rect 120862 398898 120944 399134
rect 120544 398866 120944 398898
rect 127456 399454 127696 399486
rect 127456 399218 127458 399454
rect 127694 399218 127696 399454
rect 127456 399134 127696 399218
rect 127456 398898 127458 399134
rect 127694 398898 127696 399134
rect 127456 398866 127696 398898
rect 140654 399454 140894 399486
rect 140654 399218 140656 399454
rect 140892 399218 140894 399454
rect 140654 399134 140894 399218
rect 140654 398898 140656 399134
rect 140892 398898 140894 399134
rect 140654 398866 140894 398898
rect 141500 399454 141740 399486
rect 141500 399218 141502 399454
rect 141738 399218 141740 399454
rect 141500 399134 141740 399218
rect 141500 398898 141502 399134
rect 141738 398898 141740 399134
rect 141500 398866 141740 398898
rect 147286 399454 147526 399486
rect 147286 399218 147288 399454
rect 147524 399218 147526 399454
rect 147286 399134 147526 399218
rect 147286 398898 147288 399134
rect 147524 398898 147526 399134
rect 147286 398866 147526 398898
rect 149658 399454 149898 399486
rect 149658 399218 149660 399454
rect 149896 399218 149898 399454
rect 149658 399134 149898 399218
rect 149658 398898 149660 399134
rect 149896 398898 149898 399134
rect 149658 398866 149898 398898
rect 150504 399454 150744 399486
rect 150504 399218 150506 399454
rect 150742 399218 150744 399454
rect 150504 399134 150744 399218
rect 150504 398898 150506 399134
rect 150742 398898 150744 399134
rect 150504 398866 150744 398898
rect 159504 399454 159744 399486
rect 159504 399218 159506 399454
rect 159742 399218 159744 399454
rect 159504 399134 159744 399218
rect 159504 398898 159506 399134
rect 159742 398898 159744 399134
rect 159504 398866 159744 398898
rect 168504 399454 168744 399486
rect 168504 399218 168506 399454
rect 168742 399218 168744 399454
rect 168504 399134 168744 399218
rect 168504 398898 168506 399134
rect 168742 398898 168744 399134
rect 168504 398866 168744 398898
rect 177504 399454 177744 399486
rect 177504 399218 177506 399454
rect 177742 399218 177744 399454
rect 177504 399134 177744 399218
rect 177504 398898 177506 399134
rect 177742 398898 177744 399134
rect 177504 398866 177744 398898
rect 186504 399454 186744 399486
rect 186504 399218 186506 399454
rect 186742 399218 186744 399454
rect 186504 399134 186744 399218
rect 186504 398898 186506 399134
rect 186742 398898 186744 399134
rect 186504 398866 186744 398898
rect 188306 399454 188546 399486
rect 188306 399218 188308 399454
rect 188544 399218 188546 399454
rect 188306 399134 188546 399218
rect 188306 398898 188308 399134
rect 188544 398898 188546 399134
rect 188306 398866 188546 398898
rect 190678 399454 190918 399486
rect 190678 399218 190680 399454
rect 190916 399218 190918 399454
rect 190678 399134 190918 399218
rect 190678 398898 190680 399134
rect 190916 398898 190918 399134
rect 190678 398866 190918 398898
rect 191524 399454 191764 399486
rect 191524 399218 191526 399454
rect 191762 399218 191764 399454
rect 191524 399134 191764 399218
rect 191524 398898 191526 399134
rect 191762 398898 191764 399134
rect 191524 398866 191764 398898
rect 200524 399454 200764 399486
rect 200524 399218 200526 399454
rect 200762 399218 200764 399454
rect 200524 399134 200764 399218
rect 200524 398898 200526 399134
rect 200762 398898 200764 399134
rect 200524 398866 200764 398898
rect 209524 399454 209764 399486
rect 209524 399218 209526 399454
rect 209762 399218 209764 399454
rect 209524 399134 209764 399218
rect 209524 398898 209526 399134
rect 209762 398898 209764 399134
rect 209524 398866 209764 398898
rect 218524 399454 218764 399486
rect 218524 399218 218526 399454
rect 218762 399218 218764 399454
rect 218524 399134 218764 399218
rect 218524 398898 218526 399134
rect 218762 398898 218764 399134
rect 218524 398866 218764 398898
rect 227524 399454 227764 399486
rect 227524 399218 227526 399454
rect 227762 399218 227764 399454
rect 227524 399134 227764 399218
rect 227524 398898 227526 399134
rect 227762 398898 227764 399134
rect 227524 398866 227764 398898
rect 229326 399454 229566 399486
rect 229326 399218 229328 399454
rect 229564 399218 229566 399454
rect 229326 399134 229566 399218
rect 229326 398898 229328 399134
rect 229564 398898 229566 399134
rect 229326 398866 229566 398898
rect 230698 399454 230938 399486
rect 230698 399218 230700 399454
rect 230936 399218 230938 399454
rect 230698 399134 230938 399218
rect 230698 398898 230700 399134
rect 230936 398898 230938 399134
rect 230698 398866 230938 398898
rect 231544 399454 231784 399486
rect 231544 399218 231546 399454
rect 231782 399218 231784 399454
rect 231544 399134 231784 399218
rect 231544 398898 231546 399134
rect 231782 398898 231784 399134
rect 231544 398866 231784 398898
rect 240544 399454 240784 399486
rect 240544 399218 240546 399454
rect 240782 399218 240784 399454
rect 240544 399134 240784 399218
rect 240544 398898 240546 399134
rect 240782 398898 240784 399134
rect 240544 398866 240784 398898
rect 249544 399454 249784 399486
rect 249544 399218 249546 399454
rect 249782 399218 249784 399454
rect 249544 399134 249784 399218
rect 249544 398898 249546 399134
rect 249782 398898 249784 399134
rect 249544 398866 249784 398898
rect 258544 399454 258784 399486
rect 258544 399218 258546 399454
rect 258782 399218 258784 399454
rect 258544 399134 258784 399218
rect 258544 398898 258546 399134
rect 258782 398898 258784 399134
rect 258544 398866 258784 398898
rect 267544 399454 267784 399486
rect 267544 399218 267546 399454
rect 267782 399218 267784 399454
rect 267544 399134 267784 399218
rect 267544 398898 267546 399134
rect 267782 398898 267784 399134
rect 267544 398866 267784 398898
rect 269346 399454 269586 399486
rect 269346 399218 269348 399454
rect 269584 399218 269586 399454
rect 269346 399134 269586 399218
rect 269346 398898 269348 399134
rect 269584 398898 269586 399134
rect 269346 398866 269586 398898
rect 270718 399454 270958 399486
rect 270718 399218 270720 399454
rect 270956 399218 270958 399454
rect 270718 399134 270958 399218
rect 270718 398898 270720 399134
rect 270956 398898 270958 399134
rect 270718 398866 270958 398898
rect 271564 399454 271804 399486
rect 271564 399218 271566 399454
rect 271802 399218 271804 399454
rect 271564 399134 271804 399218
rect 271564 398898 271566 399134
rect 271802 398898 271804 399134
rect 271564 398866 271804 398898
rect 280564 399454 280804 399486
rect 280564 399218 280566 399454
rect 280802 399218 280804 399454
rect 280564 399134 280804 399218
rect 280564 398898 280566 399134
rect 280802 398898 280804 399134
rect 280564 398866 280804 398898
rect 289564 399454 289804 399486
rect 289564 399218 289566 399454
rect 289802 399218 289804 399454
rect 289564 399134 289804 399218
rect 289564 398898 289566 399134
rect 289802 398898 289804 399134
rect 289564 398866 289804 398898
rect 298564 399454 298804 399486
rect 298564 399218 298566 399454
rect 298802 399218 298804 399454
rect 298564 399134 298804 399218
rect 298564 398898 298566 399134
rect 298802 398898 298804 399134
rect 298564 398866 298804 398898
rect 307564 399454 307804 399486
rect 307564 399218 307566 399454
rect 307802 399218 307804 399454
rect 307564 399134 307804 399218
rect 307564 398898 307566 399134
rect 307802 398898 307804 399134
rect 307564 398866 307804 398898
rect 309366 399454 309606 399486
rect 309366 399218 309368 399454
rect 309604 399218 309606 399454
rect 309366 399134 309606 399218
rect 309366 398898 309368 399134
rect 309604 398898 309606 399134
rect 309366 398866 309606 398898
rect 311738 399454 311978 399486
rect 311738 399218 311740 399454
rect 311976 399218 311978 399454
rect 311738 399134 311978 399218
rect 311738 398898 311740 399134
rect 311976 398898 311978 399134
rect 311738 398866 311978 398898
rect 312584 399454 312824 399486
rect 312584 399218 312586 399454
rect 312822 399218 312824 399454
rect 312584 399134 312824 399218
rect 312584 398898 312586 399134
rect 312822 398898 312824 399134
rect 312584 398866 312824 398898
rect 321584 399454 321824 399486
rect 321584 399218 321586 399454
rect 321822 399218 321824 399454
rect 321584 399134 321824 399218
rect 321584 398898 321586 399134
rect 321822 398898 321824 399134
rect 321584 398866 321824 398898
rect 330584 399454 330824 399486
rect 330584 399218 330586 399454
rect 330822 399218 330824 399454
rect 330584 399134 330824 399218
rect 330584 398898 330586 399134
rect 330822 398898 330824 399134
rect 330584 398866 330824 398898
rect 339584 399454 339824 399486
rect 339584 399218 339586 399454
rect 339822 399218 339824 399454
rect 339584 399134 339824 399218
rect 339584 398898 339586 399134
rect 339822 398898 339824 399134
rect 339584 398866 339824 398898
rect 348584 399454 348824 399486
rect 348584 399218 348586 399454
rect 348822 399218 348824 399454
rect 348584 399134 348824 399218
rect 348584 398898 348586 399134
rect 348822 398898 348824 399134
rect 348584 398866 348824 398898
rect 350386 399454 350626 399486
rect 350386 399218 350388 399454
rect 350624 399218 350626 399454
rect 350386 399134 350626 399218
rect 350386 398898 350388 399134
rect 350624 398898 350626 399134
rect 350386 398866 350626 398898
rect 352758 399454 352998 399486
rect 352758 399218 352760 399454
rect 352996 399218 352998 399454
rect 352758 399134 352998 399218
rect 352758 398898 352760 399134
rect 352996 398898 352998 399134
rect 352758 398866 352998 398898
rect 353604 399454 353844 399486
rect 353604 399218 353606 399454
rect 353842 399218 353844 399454
rect 353604 399134 353844 399218
rect 353604 398898 353606 399134
rect 353842 398898 353844 399134
rect 353604 398866 353844 398898
rect 362604 399454 362844 399486
rect 362604 399218 362606 399454
rect 362842 399218 362844 399454
rect 362604 399134 362844 399218
rect 362604 398898 362606 399134
rect 362842 398898 362844 399134
rect 362604 398866 362844 398898
rect 371604 399454 371844 399486
rect 371604 399218 371606 399454
rect 371842 399218 371844 399454
rect 371604 399134 371844 399218
rect 371604 398898 371606 399134
rect 371842 398898 371844 399134
rect 371604 398866 371844 398898
rect 380604 399454 380844 399486
rect 380604 399218 380606 399454
rect 380842 399218 380844 399454
rect 380604 399134 380844 399218
rect 380604 398898 380606 399134
rect 380842 398898 380844 399134
rect 380604 398866 380844 398898
rect 389604 399454 389844 399486
rect 389604 399218 389606 399454
rect 389842 399218 389844 399454
rect 389604 399134 389844 399218
rect 389604 398898 389606 399134
rect 389842 398898 389844 399134
rect 389604 398866 389844 398898
rect 391406 399454 391646 399486
rect 391406 399218 391408 399454
rect 391644 399218 391646 399454
rect 391406 399134 391646 399218
rect 391406 398898 391408 399134
rect 391644 398898 391646 399134
rect 391406 398866 391646 398898
rect 392778 399454 393018 399486
rect 392778 399218 392780 399454
rect 393016 399218 393018 399454
rect 392778 399134 393018 399218
rect 392778 398898 392780 399134
rect 393016 398898 393018 399134
rect 392778 398866 393018 398898
rect 393624 399454 393864 399486
rect 393624 399218 393626 399454
rect 393862 399218 393864 399454
rect 393624 399134 393864 399218
rect 393624 398898 393626 399134
rect 393862 398898 393864 399134
rect 393624 398866 393864 398898
rect 402624 399454 402864 399486
rect 402624 399218 402626 399454
rect 402862 399218 402864 399454
rect 402624 399134 402864 399218
rect 402624 398898 402626 399134
rect 402862 398898 402864 399134
rect 402624 398866 402864 398898
rect 411624 399454 411864 399486
rect 411624 399218 411626 399454
rect 411862 399218 411864 399454
rect 411624 399134 411864 399218
rect 411624 398898 411626 399134
rect 411862 398898 411864 399134
rect 411624 398866 411864 398898
rect 420624 399454 420864 399486
rect 420624 399218 420626 399454
rect 420862 399218 420864 399454
rect 420624 399134 420864 399218
rect 420624 398898 420626 399134
rect 420862 398898 420864 399134
rect 420624 398866 420864 398898
rect 429624 399454 429864 399486
rect 429624 399218 429626 399454
rect 429862 399218 429864 399454
rect 429624 399134 429864 399218
rect 429624 398898 429626 399134
rect 429862 398898 429864 399134
rect 429624 398866 429864 398898
rect 431426 399454 431666 399486
rect 431426 399218 431428 399454
rect 431664 399218 431666 399454
rect 431426 399134 431666 399218
rect 431426 398898 431428 399134
rect 431664 398898 431666 399134
rect 431426 398866 431666 398898
rect 432798 399454 433038 399486
rect 432798 399218 432800 399454
rect 433036 399218 433038 399454
rect 432798 399134 433038 399218
rect 432798 398898 432800 399134
rect 433036 398898 433038 399134
rect 432798 398866 433038 398898
rect 433644 399454 433884 399486
rect 433644 399218 433646 399454
rect 433882 399218 433884 399454
rect 433644 399134 433884 399218
rect 433644 398898 433646 399134
rect 433882 398898 433884 399134
rect 433644 398866 433884 398898
rect 439430 399454 439670 399486
rect 439430 399218 439432 399454
rect 439668 399218 439670 399454
rect 439430 399134 439670 399218
rect 439430 398898 439432 399134
rect 439668 398898 439670 399134
rect 439430 398866 439670 398898
rect 456608 399454 456848 399486
rect 456608 399218 456610 399454
rect 456846 399218 456848 399454
rect 456608 399134 456848 399218
rect 456608 398898 456610 399134
rect 456846 398898 456848 399134
rect 456608 398866 456848 398898
rect 463360 399454 463760 399486
rect 463360 399218 463442 399454
rect 463678 399218 463760 399454
rect 463360 399134 463760 399218
rect 463360 398898 463442 399134
rect 463678 398898 463760 399134
rect 463360 398866 463760 398898
rect 470648 399454 470884 399486
rect 470648 399134 470884 399218
rect 470648 398866 470884 398898
rect 479648 399454 479884 399486
rect 479648 399134 479884 399218
rect 479648 398866 479884 398898
rect 488648 399454 488884 399486
rect 488648 399134 488884 399218
rect 488648 398866 488884 398898
rect 497648 399454 497884 399486
rect 497648 399134 497884 399218
rect 497648 398866 497884 398898
rect 506648 399454 506884 399486
rect 506648 399134 506884 399218
rect 506648 398866 506884 398898
rect 515648 399454 515884 399486
rect 515648 399134 515884 399218
rect 515648 398866 515884 398898
rect 524648 399454 524884 399486
rect 524648 399134 524884 399218
rect 524648 398866 524884 398898
rect 533648 399454 533884 399486
rect 533648 399134 533884 399218
rect 533648 398866 533884 398898
rect 542648 399454 542884 399486
rect 542648 399134 542884 399218
rect 542648 398866 542884 398898
rect 551648 399454 551884 399486
rect 551648 399134 551884 399218
rect 551648 398866 551884 398898
rect 560648 399454 560884 399486
rect 560648 399134 560884 399218
rect 560648 398866 560884 398898
rect 569648 399454 569884 399486
rect 569648 399134 569884 399218
rect 569648 398866 569884 398898
rect 570768 399454 571168 399486
rect 570768 399218 570850 399454
rect 571086 399218 571168 399454
rect 570768 399134 571168 399218
rect 570768 398898 570850 399134
rect 571086 398898 571168 399134
rect 570768 398866 571168 398898
rect 578488 399454 579088 399486
rect 578488 399218 578670 399454
rect 578906 399218 579088 399454
rect 578488 399134 579088 399218
rect 578488 398898 578670 399134
rect 578906 398898 579088 399134
rect 578488 398866 579088 398898
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 4400 381454 5000 381486
rect 4400 381218 4582 381454
rect 4818 381218 5000 381454
rect 4400 381134 5000 381218
rect 4400 380898 4582 381134
rect 4818 380898 5000 381134
rect 4400 380866 5000 380898
rect 127056 381454 127296 381486
rect 127056 381218 127058 381454
rect 127294 381218 127296 381454
rect 127056 381134 127296 381218
rect 127056 380898 127058 381134
rect 127294 380898 127296 381134
rect 127056 380866 127296 380898
rect 140294 381454 140534 381486
rect 140294 381218 140296 381454
rect 140532 381218 140534 381454
rect 140294 381134 140534 381218
rect 140294 380898 140296 381134
rect 140532 380898 140534 381134
rect 140294 380866 140534 380898
rect 141100 381454 141340 381486
rect 141100 381218 141102 381454
rect 141338 381218 141340 381454
rect 141100 381134 141340 381218
rect 141100 380898 141102 381134
rect 141338 380898 141340 381134
rect 141100 380866 141340 380898
rect 147646 381454 147886 381486
rect 147646 381218 147648 381454
rect 147884 381218 147886 381454
rect 147646 381134 147886 381218
rect 147646 380898 147648 381134
rect 147884 380898 147886 381134
rect 147646 380866 147886 380898
rect 149298 381454 149538 381486
rect 149298 381218 149300 381454
rect 149536 381218 149538 381454
rect 149298 381134 149538 381218
rect 149298 380898 149300 381134
rect 149536 380898 149538 381134
rect 149298 380866 149538 380898
rect 150104 381454 150344 381486
rect 150104 381218 150106 381454
rect 150342 381218 150344 381454
rect 150104 381134 150344 381218
rect 150104 380898 150106 381134
rect 150342 380898 150344 381134
rect 150104 380866 150344 380898
rect 159104 381454 159344 381486
rect 159104 381218 159106 381454
rect 159342 381218 159344 381454
rect 159104 381134 159344 381218
rect 159104 380898 159106 381134
rect 159342 380898 159344 381134
rect 159104 380866 159344 380898
rect 168104 381454 168344 381486
rect 168104 381218 168106 381454
rect 168342 381218 168344 381454
rect 168104 381134 168344 381218
rect 168104 380898 168106 381134
rect 168342 380898 168344 381134
rect 168104 380866 168344 380898
rect 177104 381454 177344 381486
rect 177104 381218 177106 381454
rect 177342 381218 177344 381454
rect 177104 381134 177344 381218
rect 177104 380898 177106 381134
rect 177342 380898 177344 381134
rect 177104 380866 177344 380898
rect 186104 381454 186344 381486
rect 186104 381218 186106 381454
rect 186342 381218 186344 381454
rect 186104 381134 186344 381218
rect 186104 380898 186106 381134
rect 186342 380898 186344 381134
rect 186104 380866 186344 380898
rect 188666 381454 188906 381486
rect 188666 381218 188668 381454
rect 188904 381218 188906 381454
rect 188666 381134 188906 381218
rect 188666 380898 188668 381134
rect 188904 380898 188906 381134
rect 188666 380866 188906 380898
rect 190318 381454 190558 381486
rect 190318 381218 190320 381454
rect 190556 381218 190558 381454
rect 190318 381134 190558 381218
rect 190318 380898 190320 381134
rect 190556 380898 190558 381134
rect 190318 380866 190558 380898
rect 191124 381454 191364 381486
rect 191124 381218 191126 381454
rect 191362 381218 191364 381454
rect 191124 381134 191364 381218
rect 191124 380898 191126 381134
rect 191362 380898 191364 381134
rect 191124 380866 191364 380898
rect 200124 381454 200364 381486
rect 200124 381218 200126 381454
rect 200362 381218 200364 381454
rect 200124 381134 200364 381218
rect 200124 380898 200126 381134
rect 200362 380898 200364 381134
rect 200124 380866 200364 380898
rect 209124 381454 209364 381486
rect 209124 381218 209126 381454
rect 209362 381218 209364 381454
rect 209124 381134 209364 381218
rect 209124 380898 209126 381134
rect 209362 380898 209364 381134
rect 209124 380866 209364 380898
rect 218124 381454 218364 381486
rect 218124 381218 218126 381454
rect 218362 381218 218364 381454
rect 218124 381134 218364 381218
rect 218124 380898 218126 381134
rect 218362 380898 218364 381134
rect 218124 380866 218364 380898
rect 227124 381454 227364 381486
rect 227124 381218 227126 381454
rect 227362 381218 227364 381454
rect 227124 381134 227364 381218
rect 227124 380898 227126 381134
rect 227362 380898 227364 381134
rect 227124 380866 227364 380898
rect 229686 381454 229926 381486
rect 229686 381218 229688 381454
rect 229924 381218 229926 381454
rect 229686 381134 229926 381218
rect 229686 380898 229688 381134
rect 229924 380898 229926 381134
rect 229686 380866 229926 380898
rect 230338 381454 230578 381486
rect 230338 381218 230340 381454
rect 230576 381218 230578 381454
rect 230338 381134 230578 381218
rect 230338 380898 230340 381134
rect 230576 380898 230578 381134
rect 230338 380866 230578 380898
rect 231144 381454 231384 381486
rect 231144 381218 231146 381454
rect 231382 381218 231384 381454
rect 231144 381134 231384 381218
rect 231144 380898 231146 381134
rect 231382 380898 231384 381134
rect 231144 380866 231384 380898
rect 240144 381454 240384 381486
rect 240144 381218 240146 381454
rect 240382 381218 240384 381454
rect 240144 381134 240384 381218
rect 240144 380898 240146 381134
rect 240382 380898 240384 381134
rect 240144 380866 240384 380898
rect 249144 381454 249384 381486
rect 249144 381218 249146 381454
rect 249382 381218 249384 381454
rect 249144 381134 249384 381218
rect 249144 380898 249146 381134
rect 249382 380898 249384 381134
rect 249144 380866 249384 380898
rect 258144 381454 258384 381486
rect 258144 381218 258146 381454
rect 258382 381218 258384 381454
rect 258144 381134 258384 381218
rect 258144 380898 258146 381134
rect 258382 380898 258384 381134
rect 258144 380866 258384 380898
rect 267144 381454 267384 381486
rect 267144 381218 267146 381454
rect 267382 381218 267384 381454
rect 267144 381134 267384 381218
rect 267144 380898 267146 381134
rect 267382 380898 267384 381134
rect 267144 380866 267384 380898
rect 269706 381454 269946 381486
rect 269706 381218 269708 381454
rect 269944 381218 269946 381454
rect 269706 381134 269946 381218
rect 269706 380898 269708 381134
rect 269944 380898 269946 381134
rect 269706 380866 269946 380898
rect 270358 381454 270598 381486
rect 270358 381218 270360 381454
rect 270596 381218 270598 381454
rect 270358 381134 270598 381218
rect 270358 380898 270360 381134
rect 270596 380898 270598 381134
rect 270358 380866 270598 380898
rect 271164 381454 271404 381486
rect 271164 381218 271166 381454
rect 271402 381218 271404 381454
rect 271164 381134 271404 381218
rect 271164 380898 271166 381134
rect 271402 380898 271404 381134
rect 271164 380866 271404 380898
rect 280164 381454 280404 381486
rect 280164 381218 280166 381454
rect 280402 381218 280404 381454
rect 280164 381134 280404 381218
rect 280164 380898 280166 381134
rect 280402 380898 280404 381134
rect 280164 380866 280404 380898
rect 289164 381454 289404 381486
rect 289164 381218 289166 381454
rect 289402 381218 289404 381454
rect 289164 381134 289404 381218
rect 289164 380898 289166 381134
rect 289402 380898 289404 381134
rect 289164 380866 289404 380898
rect 298164 381454 298404 381486
rect 298164 381218 298166 381454
rect 298402 381218 298404 381454
rect 298164 381134 298404 381218
rect 298164 380898 298166 381134
rect 298402 380898 298404 381134
rect 298164 380866 298404 380898
rect 307164 381454 307404 381486
rect 307164 381218 307166 381454
rect 307402 381218 307404 381454
rect 307164 381134 307404 381218
rect 307164 380898 307166 381134
rect 307402 380898 307404 381134
rect 307164 380866 307404 380898
rect 309726 381454 309966 381486
rect 309726 381218 309728 381454
rect 309964 381218 309966 381454
rect 309726 381134 309966 381218
rect 309726 380898 309728 381134
rect 309964 380898 309966 381134
rect 309726 380866 309966 380898
rect 311378 381454 311618 381486
rect 311378 381218 311380 381454
rect 311616 381218 311618 381454
rect 311378 381134 311618 381218
rect 311378 380898 311380 381134
rect 311616 380898 311618 381134
rect 311378 380866 311618 380898
rect 312184 381454 312424 381486
rect 312184 381218 312186 381454
rect 312422 381218 312424 381454
rect 312184 381134 312424 381218
rect 312184 380898 312186 381134
rect 312422 380898 312424 381134
rect 312184 380866 312424 380898
rect 321184 381454 321424 381486
rect 321184 381218 321186 381454
rect 321422 381218 321424 381454
rect 321184 381134 321424 381218
rect 321184 380898 321186 381134
rect 321422 380898 321424 381134
rect 321184 380866 321424 380898
rect 330184 381454 330424 381486
rect 330184 381218 330186 381454
rect 330422 381218 330424 381454
rect 330184 381134 330424 381218
rect 330184 380898 330186 381134
rect 330422 380898 330424 381134
rect 330184 380866 330424 380898
rect 339184 381454 339424 381486
rect 339184 381218 339186 381454
rect 339422 381218 339424 381454
rect 339184 381134 339424 381218
rect 339184 380898 339186 381134
rect 339422 380898 339424 381134
rect 339184 380866 339424 380898
rect 348184 381454 348424 381486
rect 348184 381218 348186 381454
rect 348422 381218 348424 381454
rect 348184 381134 348424 381218
rect 348184 380898 348186 381134
rect 348422 380898 348424 381134
rect 348184 380866 348424 380898
rect 350746 381454 350986 381486
rect 350746 381218 350748 381454
rect 350984 381218 350986 381454
rect 350746 381134 350986 381218
rect 350746 380898 350748 381134
rect 350984 380898 350986 381134
rect 350746 380866 350986 380898
rect 352398 381454 352638 381486
rect 352398 381218 352400 381454
rect 352636 381218 352638 381454
rect 352398 381134 352638 381218
rect 352398 380898 352400 381134
rect 352636 380898 352638 381134
rect 352398 380866 352638 380898
rect 353204 381454 353444 381486
rect 353204 381218 353206 381454
rect 353442 381218 353444 381454
rect 353204 381134 353444 381218
rect 353204 380898 353206 381134
rect 353442 380898 353444 381134
rect 353204 380866 353444 380898
rect 362204 381454 362444 381486
rect 362204 381218 362206 381454
rect 362442 381218 362444 381454
rect 362204 381134 362444 381218
rect 362204 380898 362206 381134
rect 362442 380898 362444 381134
rect 362204 380866 362444 380898
rect 371204 381454 371444 381486
rect 371204 381218 371206 381454
rect 371442 381218 371444 381454
rect 371204 381134 371444 381218
rect 371204 380898 371206 381134
rect 371442 380898 371444 381134
rect 371204 380866 371444 380898
rect 380204 381454 380444 381486
rect 380204 381218 380206 381454
rect 380442 381218 380444 381454
rect 380204 381134 380444 381218
rect 380204 380898 380206 381134
rect 380442 380898 380444 381134
rect 380204 380866 380444 380898
rect 389204 381454 389444 381486
rect 389204 381218 389206 381454
rect 389442 381218 389444 381454
rect 389204 381134 389444 381218
rect 389204 380898 389206 381134
rect 389442 380898 389444 381134
rect 389204 380866 389444 380898
rect 391766 381454 392006 381486
rect 391766 381218 391768 381454
rect 392004 381218 392006 381454
rect 391766 381134 392006 381218
rect 391766 380898 391768 381134
rect 392004 380898 392006 381134
rect 391766 380866 392006 380898
rect 392418 381454 392658 381486
rect 392418 381218 392420 381454
rect 392656 381218 392658 381454
rect 392418 381134 392658 381218
rect 392418 380898 392420 381134
rect 392656 380898 392658 381134
rect 392418 380866 392658 380898
rect 393224 381454 393464 381486
rect 393224 381218 393226 381454
rect 393462 381218 393464 381454
rect 393224 381134 393464 381218
rect 393224 380898 393226 381134
rect 393462 380898 393464 381134
rect 393224 380866 393464 380898
rect 402224 381454 402464 381486
rect 402224 381218 402226 381454
rect 402462 381218 402464 381454
rect 402224 381134 402464 381218
rect 402224 380898 402226 381134
rect 402462 380898 402464 381134
rect 402224 380866 402464 380898
rect 411224 381454 411464 381486
rect 411224 381218 411226 381454
rect 411462 381218 411464 381454
rect 411224 381134 411464 381218
rect 411224 380898 411226 381134
rect 411462 380898 411464 381134
rect 411224 380866 411464 380898
rect 420224 381454 420464 381486
rect 420224 381218 420226 381454
rect 420462 381218 420464 381454
rect 420224 381134 420464 381218
rect 420224 380898 420226 381134
rect 420462 380898 420464 381134
rect 420224 380866 420464 380898
rect 429224 381454 429464 381486
rect 429224 381218 429226 381454
rect 429462 381218 429464 381454
rect 429224 381134 429464 381218
rect 429224 380898 429226 381134
rect 429462 380898 429464 381134
rect 429224 380866 429464 380898
rect 431786 381454 432026 381486
rect 431786 381218 431788 381454
rect 432024 381218 432026 381454
rect 431786 381134 432026 381218
rect 431786 380898 431788 381134
rect 432024 380898 432026 381134
rect 431786 380866 432026 380898
rect 432438 381454 432678 381486
rect 432438 381218 432440 381454
rect 432676 381218 432678 381454
rect 432438 381134 432678 381218
rect 432438 380898 432440 381134
rect 432676 380898 432678 381134
rect 432438 380866 432678 380898
rect 433244 381454 433484 381486
rect 433244 381218 433246 381454
rect 433482 381218 433484 381454
rect 433244 381134 433484 381218
rect 433244 380898 433246 381134
rect 433482 380898 433484 381134
rect 433244 380866 433484 380898
rect 439790 381454 440030 381486
rect 439790 381218 439792 381454
rect 440028 381218 440030 381454
rect 439790 381134 440030 381218
rect 439790 380898 439792 381134
rect 440028 380898 440030 381134
rect 439790 380866 440030 380898
rect 457008 381454 457248 381486
rect 457008 381218 457010 381454
rect 457246 381218 457248 381454
rect 457008 381134 457248 381218
rect 457008 380898 457010 381134
rect 457246 380898 457248 381134
rect 457008 380866 457248 380898
rect 579288 381454 579888 381486
rect 579288 381218 579470 381454
rect 579706 381218 579888 381454
rect 579288 381134 579888 381218
rect 579288 380898 579470 381134
rect 579706 380898 579888 381134
rect 579288 380866 579888 380898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect 5200 363454 5800 363486
rect 5200 363218 5382 363454
rect 5618 363218 5800 363454
rect 5200 363134 5800 363218
rect 5200 362898 5382 363134
rect 5618 362898 5800 363134
rect 5200 362866 5800 362898
rect 127456 363454 127696 363486
rect 127456 363218 127458 363454
rect 127694 363218 127696 363454
rect 127456 363134 127696 363218
rect 127456 362898 127458 363134
rect 127694 362898 127696 363134
rect 127456 362866 127696 362898
rect 140654 363454 140894 363486
rect 140654 363218 140656 363454
rect 140892 363218 140894 363454
rect 140654 363134 140894 363218
rect 140654 362898 140656 363134
rect 140892 362898 140894 363134
rect 140654 362866 140894 362898
rect 141500 363454 141740 363486
rect 141500 363218 141502 363454
rect 141738 363218 141740 363454
rect 141500 363134 141740 363218
rect 141500 362898 141502 363134
rect 141738 362898 141740 363134
rect 141500 362866 141740 362898
rect 147286 363454 147526 363486
rect 147286 363218 147288 363454
rect 147524 363218 147526 363454
rect 147286 363134 147526 363218
rect 147286 362898 147288 363134
rect 147524 362898 147526 363134
rect 147286 362866 147526 362898
rect 149658 363454 149898 363486
rect 149658 363218 149660 363454
rect 149896 363218 149898 363454
rect 149658 363134 149898 363218
rect 149658 362898 149660 363134
rect 149896 362898 149898 363134
rect 149658 362866 149898 362898
rect 150504 363454 150744 363486
rect 150504 363218 150506 363454
rect 150742 363218 150744 363454
rect 150504 363134 150744 363218
rect 150504 362898 150506 363134
rect 150742 362898 150744 363134
rect 150504 362866 150744 362898
rect 159504 363454 159744 363486
rect 159504 363218 159506 363454
rect 159742 363218 159744 363454
rect 159504 363134 159744 363218
rect 159504 362898 159506 363134
rect 159742 362898 159744 363134
rect 159504 362866 159744 362898
rect 168504 363454 168744 363486
rect 168504 363218 168506 363454
rect 168742 363218 168744 363454
rect 168504 363134 168744 363218
rect 168504 362898 168506 363134
rect 168742 362898 168744 363134
rect 168504 362866 168744 362898
rect 177504 363454 177744 363486
rect 177504 363218 177506 363454
rect 177742 363218 177744 363454
rect 177504 363134 177744 363218
rect 177504 362898 177506 363134
rect 177742 362898 177744 363134
rect 177504 362866 177744 362898
rect 186504 363454 186744 363486
rect 186504 363218 186506 363454
rect 186742 363218 186744 363454
rect 186504 363134 186744 363218
rect 186504 362898 186506 363134
rect 186742 362898 186744 363134
rect 186504 362866 186744 362898
rect 188306 363454 188546 363486
rect 188306 363218 188308 363454
rect 188544 363218 188546 363454
rect 188306 363134 188546 363218
rect 188306 362898 188308 363134
rect 188544 362898 188546 363134
rect 188306 362866 188546 362898
rect 190678 363454 190918 363486
rect 190678 363218 190680 363454
rect 190916 363218 190918 363454
rect 190678 363134 190918 363218
rect 190678 362898 190680 363134
rect 190916 362898 190918 363134
rect 190678 362866 190918 362898
rect 191524 363454 191764 363486
rect 191524 363218 191526 363454
rect 191762 363218 191764 363454
rect 191524 363134 191764 363218
rect 191524 362898 191526 363134
rect 191762 362898 191764 363134
rect 191524 362866 191764 362898
rect 200524 363454 200764 363486
rect 200524 363218 200526 363454
rect 200762 363218 200764 363454
rect 200524 363134 200764 363218
rect 200524 362898 200526 363134
rect 200762 362898 200764 363134
rect 200524 362866 200764 362898
rect 209524 363454 209764 363486
rect 209524 363218 209526 363454
rect 209762 363218 209764 363454
rect 209524 363134 209764 363218
rect 209524 362898 209526 363134
rect 209762 362898 209764 363134
rect 209524 362866 209764 362898
rect 218524 363454 218764 363486
rect 218524 363218 218526 363454
rect 218762 363218 218764 363454
rect 218524 363134 218764 363218
rect 218524 362898 218526 363134
rect 218762 362898 218764 363134
rect 218524 362866 218764 362898
rect 227524 363454 227764 363486
rect 227524 363218 227526 363454
rect 227762 363218 227764 363454
rect 227524 363134 227764 363218
rect 227524 362898 227526 363134
rect 227762 362898 227764 363134
rect 227524 362866 227764 362898
rect 229326 363454 229566 363486
rect 229326 363218 229328 363454
rect 229564 363218 229566 363454
rect 229326 363134 229566 363218
rect 229326 362898 229328 363134
rect 229564 362898 229566 363134
rect 229326 362866 229566 362898
rect 230698 363454 230938 363486
rect 230698 363218 230700 363454
rect 230936 363218 230938 363454
rect 230698 363134 230938 363218
rect 230698 362898 230700 363134
rect 230936 362898 230938 363134
rect 230698 362866 230938 362898
rect 231544 363454 231784 363486
rect 231544 363218 231546 363454
rect 231782 363218 231784 363454
rect 231544 363134 231784 363218
rect 231544 362898 231546 363134
rect 231782 362898 231784 363134
rect 231544 362866 231784 362898
rect 240544 363454 240784 363486
rect 240544 363218 240546 363454
rect 240782 363218 240784 363454
rect 240544 363134 240784 363218
rect 240544 362898 240546 363134
rect 240782 362898 240784 363134
rect 240544 362866 240784 362898
rect 249544 363454 249784 363486
rect 249544 363218 249546 363454
rect 249782 363218 249784 363454
rect 249544 363134 249784 363218
rect 249544 362898 249546 363134
rect 249782 362898 249784 363134
rect 249544 362866 249784 362898
rect 258544 363454 258784 363486
rect 258544 363218 258546 363454
rect 258782 363218 258784 363454
rect 258544 363134 258784 363218
rect 258544 362898 258546 363134
rect 258782 362898 258784 363134
rect 258544 362866 258784 362898
rect 267544 363454 267784 363486
rect 267544 363218 267546 363454
rect 267782 363218 267784 363454
rect 267544 363134 267784 363218
rect 267544 362898 267546 363134
rect 267782 362898 267784 363134
rect 267544 362866 267784 362898
rect 269346 363454 269586 363486
rect 269346 363218 269348 363454
rect 269584 363218 269586 363454
rect 269346 363134 269586 363218
rect 269346 362898 269348 363134
rect 269584 362898 269586 363134
rect 269346 362866 269586 362898
rect 270718 363454 270958 363486
rect 270718 363218 270720 363454
rect 270956 363218 270958 363454
rect 270718 363134 270958 363218
rect 270718 362898 270720 363134
rect 270956 362898 270958 363134
rect 270718 362866 270958 362898
rect 271564 363454 271804 363486
rect 271564 363218 271566 363454
rect 271802 363218 271804 363454
rect 271564 363134 271804 363218
rect 271564 362898 271566 363134
rect 271802 362898 271804 363134
rect 271564 362866 271804 362898
rect 280564 363454 280804 363486
rect 280564 363218 280566 363454
rect 280802 363218 280804 363454
rect 280564 363134 280804 363218
rect 280564 362898 280566 363134
rect 280802 362898 280804 363134
rect 280564 362866 280804 362898
rect 289564 363454 289804 363486
rect 289564 363218 289566 363454
rect 289802 363218 289804 363454
rect 289564 363134 289804 363218
rect 289564 362898 289566 363134
rect 289802 362898 289804 363134
rect 289564 362866 289804 362898
rect 298564 363454 298804 363486
rect 298564 363218 298566 363454
rect 298802 363218 298804 363454
rect 298564 363134 298804 363218
rect 298564 362898 298566 363134
rect 298802 362898 298804 363134
rect 298564 362866 298804 362898
rect 307564 363454 307804 363486
rect 307564 363218 307566 363454
rect 307802 363218 307804 363454
rect 307564 363134 307804 363218
rect 307564 362898 307566 363134
rect 307802 362898 307804 363134
rect 307564 362866 307804 362898
rect 309366 363454 309606 363486
rect 309366 363218 309368 363454
rect 309604 363218 309606 363454
rect 309366 363134 309606 363218
rect 309366 362898 309368 363134
rect 309604 362898 309606 363134
rect 309366 362866 309606 362898
rect 311738 363454 311978 363486
rect 311738 363218 311740 363454
rect 311976 363218 311978 363454
rect 311738 363134 311978 363218
rect 311738 362898 311740 363134
rect 311976 362898 311978 363134
rect 311738 362866 311978 362898
rect 312584 363454 312824 363486
rect 312584 363218 312586 363454
rect 312822 363218 312824 363454
rect 312584 363134 312824 363218
rect 312584 362898 312586 363134
rect 312822 362898 312824 363134
rect 312584 362866 312824 362898
rect 321584 363454 321824 363486
rect 321584 363218 321586 363454
rect 321822 363218 321824 363454
rect 321584 363134 321824 363218
rect 321584 362898 321586 363134
rect 321822 362898 321824 363134
rect 321584 362866 321824 362898
rect 330584 363454 330824 363486
rect 330584 363218 330586 363454
rect 330822 363218 330824 363454
rect 330584 363134 330824 363218
rect 330584 362898 330586 363134
rect 330822 362898 330824 363134
rect 330584 362866 330824 362898
rect 339584 363454 339824 363486
rect 339584 363218 339586 363454
rect 339822 363218 339824 363454
rect 339584 363134 339824 363218
rect 339584 362898 339586 363134
rect 339822 362898 339824 363134
rect 339584 362866 339824 362898
rect 348584 363454 348824 363486
rect 348584 363218 348586 363454
rect 348822 363218 348824 363454
rect 348584 363134 348824 363218
rect 348584 362898 348586 363134
rect 348822 362898 348824 363134
rect 348584 362866 348824 362898
rect 350386 363454 350626 363486
rect 350386 363218 350388 363454
rect 350624 363218 350626 363454
rect 350386 363134 350626 363218
rect 350386 362898 350388 363134
rect 350624 362898 350626 363134
rect 350386 362866 350626 362898
rect 352758 363454 352998 363486
rect 352758 363218 352760 363454
rect 352996 363218 352998 363454
rect 352758 363134 352998 363218
rect 352758 362898 352760 363134
rect 352996 362898 352998 363134
rect 352758 362866 352998 362898
rect 353604 363454 353844 363486
rect 353604 363218 353606 363454
rect 353842 363218 353844 363454
rect 353604 363134 353844 363218
rect 353604 362898 353606 363134
rect 353842 362898 353844 363134
rect 353604 362866 353844 362898
rect 362604 363454 362844 363486
rect 362604 363218 362606 363454
rect 362842 363218 362844 363454
rect 362604 363134 362844 363218
rect 362604 362898 362606 363134
rect 362842 362898 362844 363134
rect 362604 362866 362844 362898
rect 371604 363454 371844 363486
rect 371604 363218 371606 363454
rect 371842 363218 371844 363454
rect 371604 363134 371844 363218
rect 371604 362898 371606 363134
rect 371842 362898 371844 363134
rect 371604 362866 371844 362898
rect 380604 363454 380844 363486
rect 380604 363218 380606 363454
rect 380842 363218 380844 363454
rect 380604 363134 380844 363218
rect 380604 362898 380606 363134
rect 380842 362898 380844 363134
rect 380604 362866 380844 362898
rect 389604 363454 389844 363486
rect 389604 363218 389606 363454
rect 389842 363218 389844 363454
rect 389604 363134 389844 363218
rect 389604 362898 389606 363134
rect 389842 362898 389844 363134
rect 389604 362866 389844 362898
rect 391406 363454 391646 363486
rect 391406 363218 391408 363454
rect 391644 363218 391646 363454
rect 391406 363134 391646 363218
rect 391406 362898 391408 363134
rect 391644 362898 391646 363134
rect 391406 362866 391646 362898
rect 392778 363454 393018 363486
rect 392778 363218 392780 363454
rect 393016 363218 393018 363454
rect 392778 363134 393018 363218
rect 392778 362898 392780 363134
rect 393016 362898 393018 363134
rect 392778 362866 393018 362898
rect 393624 363454 393864 363486
rect 393624 363218 393626 363454
rect 393862 363218 393864 363454
rect 393624 363134 393864 363218
rect 393624 362898 393626 363134
rect 393862 362898 393864 363134
rect 393624 362866 393864 362898
rect 402624 363454 402864 363486
rect 402624 363218 402626 363454
rect 402862 363218 402864 363454
rect 402624 363134 402864 363218
rect 402624 362898 402626 363134
rect 402862 362898 402864 363134
rect 402624 362866 402864 362898
rect 411624 363454 411864 363486
rect 411624 363218 411626 363454
rect 411862 363218 411864 363454
rect 411624 363134 411864 363218
rect 411624 362898 411626 363134
rect 411862 362898 411864 363134
rect 411624 362866 411864 362898
rect 420624 363454 420864 363486
rect 420624 363218 420626 363454
rect 420862 363218 420864 363454
rect 420624 363134 420864 363218
rect 420624 362898 420626 363134
rect 420862 362898 420864 363134
rect 420624 362866 420864 362898
rect 429624 363454 429864 363486
rect 429624 363218 429626 363454
rect 429862 363218 429864 363454
rect 429624 363134 429864 363218
rect 429624 362898 429626 363134
rect 429862 362898 429864 363134
rect 429624 362866 429864 362898
rect 431426 363454 431666 363486
rect 431426 363218 431428 363454
rect 431664 363218 431666 363454
rect 431426 363134 431666 363218
rect 431426 362898 431428 363134
rect 431664 362898 431666 363134
rect 431426 362866 431666 362898
rect 432798 363454 433038 363486
rect 432798 363218 432800 363454
rect 433036 363218 433038 363454
rect 432798 363134 433038 363218
rect 432798 362898 432800 363134
rect 433036 362898 433038 363134
rect 432798 362866 433038 362898
rect 433644 363454 433884 363486
rect 433644 363218 433646 363454
rect 433882 363218 433884 363454
rect 433644 363134 433884 363218
rect 433644 362898 433646 363134
rect 433882 362898 433884 363134
rect 433644 362866 433884 362898
rect 439430 363454 439670 363486
rect 439430 363218 439432 363454
rect 439668 363218 439670 363454
rect 439430 363134 439670 363218
rect 439430 362898 439432 363134
rect 439668 362898 439670 363134
rect 439430 362866 439670 362898
rect 456608 363454 456848 363486
rect 456608 363218 456610 363454
rect 456846 363218 456848 363454
rect 456608 363134 456848 363218
rect 456608 362898 456610 363134
rect 456846 362898 456848 363134
rect 456608 362866 456848 362898
rect 578488 363454 579088 363486
rect 578488 363218 578670 363454
rect 578906 363218 579088 363454
rect 578488 363134 579088 363218
rect 578488 362898 578670 363134
rect 578906 362898 579088 363134
rect 578488 362866 579088 362898
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 4400 345454 5000 345486
rect 4400 345218 4582 345454
rect 4818 345218 5000 345454
rect 4400 345134 5000 345218
rect 4400 344898 4582 345134
rect 4818 344898 5000 345134
rect 4400 344866 5000 344898
rect 127056 345454 127296 345486
rect 127056 345218 127058 345454
rect 127294 345218 127296 345454
rect 127056 345134 127296 345218
rect 127056 344898 127058 345134
rect 127294 344898 127296 345134
rect 127056 344866 127296 344898
rect 140294 345454 140534 345486
rect 140294 345218 140296 345454
rect 140532 345218 140534 345454
rect 140294 345134 140534 345218
rect 140294 344898 140296 345134
rect 140532 344898 140534 345134
rect 140294 344866 140534 344898
rect 141100 345454 141340 345486
rect 141100 345218 141102 345454
rect 141338 345218 141340 345454
rect 141100 345134 141340 345218
rect 141100 344898 141102 345134
rect 141338 344898 141340 345134
rect 141100 344866 141340 344898
rect 147646 345454 147886 345486
rect 147646 345218 147648 345454
rect 147884 345218 147886 345454
rect 147646 345134 147886 345218
rect 147646 344898 147648 345134
rect 147884 344898 147886 345134
rect 147646 344866 147886 344898
rect 149298 345454 149538 345486
rect 149298 345218 149300 345454
rect 149536 345218 149538 345454
rect 149298 345134 149538 345218
rect 149298 344898 149300 345134
rect 149536 344898 149538 345134
rect 149298 344866 149538 344898
rect 150104 345454 150344 345486
rect 150104 345218 150106 345454
rect 150342 345218 150344 345454
rect 150104 345134 150344 345218
rect 150104 344898 150106 345134
rect 150342 344898 150344 345134
rect 150104 344866 150344 344898
rect 159104 345454 159344 345486
rect 159104 345218 159106 345454
rect 159342 345218 159344 345454
rect 159104 345134 159344 345218
rect 159104 344898 159106 345134
rect 159342 344898 159344 345134
rect 159104 344866 159344 344898
rect 168104 345454 168344 345486
rect 168104 345218 168106 345454
rect 168342 345218 168344 345454
rect 168104 345134 168344 345218
rect 168104 344898 168106 345134
rect 168342 344898 168344 345134
rect 168104 344866 168344 344898
rect 177104 345454 177344 345486
rect 177104 345218 177106 345454
rect 177342 345218 177344 345454
rect 177104 345134 177344 345218
rect 177104 344898 177106 345134
rect 177342 344898 177344 345134
rect 177104 344866 177344 344898
rect 186104 345454 186344 345486
rect 186104 345218 186106 345454
rect 186342 345218 186344 345454
rect 186104 345134 186344 345218
rect 186104 344898 186106 345134
rect 186342 344898 186344 345134
rect 186104 344866 186344 344898
rect 188666 345454 188906 345486
rect 188666 345218 188668 345454
rect 188904 345218 188906 345454
rect 188666 345134 188906 345218
rect 188666 344898 188668 345134
rect 188904 344898 188906 345134
rect 188666 344866 188906 344898
rect 190318 345454 190558 345486
rect 190318 345218 190320 345454
rect 190556 345218 190558 345454
rect 190318 345134 190558 345218
rect 190318 344898 190320 345134
rect 190556 344898 190558 345134
rect 190318 344866 190558 344898
rect 191124 345454 191364 345486
rect 191124 345218 191126 345454
rect 191362 345218 191364 345454
rect 191124 345134 191364 345218
rect 191124 344898 191126 345134
rect 191362 344898 191364 345134
rect 191124 344866 191364 344898
rect 200124 345454 200364 345486
rect 200124 345218 200126 345454
rect 200362 345218 200364 345454
rect 200124 345134 200364 345218
rect 200124 344898 200126 345134
rect 200362 344898 200364 345134
rect 200124 344866 200364 344898
rect 209124 345454 209364 345486
rect 209124 345218 209126 345454
rect 209362 345218 209364 345454
rect 209124 345134 209364 345218
rect 209124 344898 209126 345134
rect 209362 344898 209364 345134
rect 209124 344866 209364 344898
rect 218124 345454 218364 345486
rect 218124 345218 218126 345454
rect 218362 345218 218364 345454
rect 218124 345134 218364 345218
rect 218124 344898 218126 345134
rect 218362 344898 218364 345134
rect 218124 344866 218364 344898
rect 227124 345454 227364 345486
rect 227124 345218 227126 345454
rect 227362 345218 227364 345454
rect 227124 345134 227364 345218
rect 227124 344898 227126 345134
rect 227362 344898 227364 345134
rect 227124 344866 227364 344898
rect 229686 345454 229926 345486
rect 229686 345218 229688 345454
rect 229924 345218 229926 345454
rect 229686 345134 229926 345218
rect 229686 344898 229688 345134
rect 229924 344898 229926 345134
rect 229686 344866 229926 344898
rect 230338 345454 230578 345486
rect 230338 345218 230340 345454
rect 230576 345218 230578 345454
rect 230338 345134 230578 345218
rect 230338 344898 230340 345134
rect 230576 344898 230578 345134
rect 230338 344866 230578 344898
rect 231144 345454 231384 345486
rect 231144 345218 231146 345454
rect 231382 345218 231384 345454
rect 231144 345134 231384 345218
rect 231144 344898 231146 345134
rect 231382 344898 231384 345134
rect 231144 344866 231384 344898
rect 240144 345454 240384 345486
rect 240144 345218 240146 345454
rect 240382 345218 240384 345454
rect 240144 345134 240384 345218
rect 240144 344898 240146 345134
rect 240382 344898 240384 345134
rect 240144 344866 240384 344898
rect 249144 345454 249384 345486
rect 249144 345218 249146 345454
rect 249382 345218 249384 345454
rect 249144 345134 249384 345218
rect 249144 344898 249146 345134
rect 249382 344898 249384 345134
rect 249144 344866 249384 344898
rect 258144 345454 258384 345486
rect 258144 345218 258146 345454
rect 258382 345218 258384 345454
rect 258144 345134 258384 345218
rect 258144 344898 258146 345134
rect 258382 344898 258384 345134
rect 258144 344866 258384 344898
rect 267144 345454 267384 345486
rect 267144 345218 267146 345454
rect 267382 345218 267384 345454
rect 267144 345134 267384 345218
rect 267144 344898 267146 345134
rect 267382 344898 267384 345134
rect 267144 344866 267384 344898
rect 269706 345454 269946 345486
rect 269706 345218 269708 345454
rect 269944 345218 269946 345454
rect 269706 345134 269946 345218
rect 269706 344898 269708 345134
rect 269944 344898 269946 345134
rect 269706 344866 269946 344898
rect 270358 345454 270598 345486
rect 270358 345218 270360 345454
rect 270596 345218 270598 345454
rect 270358 345134 270598 345218
rect 270358 344898 270360 345134
rect 270596 344898 270598 345134
rect 270358 344866 270598 344898
rect 271164 345454 271404 345486
rect 271164 345218 271166 345454
rect 271402 345218 271404 345454
rect 271164 345134 271404 345218
rect 271164 344898 271166 345134
rect 271402 344898 271404 345134
rect 271164 344866 271404 344898
rect 280164 345454 280404 345486
rect 280164 345218 280166 345454
rect 280402 345218 280404 345454
rect 280164 345134 280404 345218
rect 280164 344898 280166 345134
rect 280402 344898 280404 345134
rect 280164 344866 280404 344898
rect 289164 345454 289404 345486
rect 289164 345218 289166 345454
rect 289402 345218 289404 345454
rect 289164 345134 289404 345218
rect 289164 344898 289166 345134
rect 289402 344898 289404 345134
rect 289164 344866 289404 344898
rect 298164 345454 298404 345486
rect 298164 345218 298166 345454
rect 298402 345218 298404 345454
rect 298164 345134 298404 345218
rect 298164 344898 298166 345134
rect 298402 344898 298404 345134
rect 298164 344866 298404 344898
rect 307164 345454 307404 345486
rect 307164 345218 307166 345454
rect 307402 345218 307404 345454
rect 307164 345134 307404 345218
rect 307164 344898 307166 345134
rect 307402 344898 307404 345134
rect 307164 344866 307404 344898
rect 309726 345454 309966 345486
rect 309726 345218 309728 345454
rect 309964 345218 309966 345454
rect 309726 345134 309966 345218
rect 309726 344898 309728 345134
rect 309964 344898 309966 345134
rect 309726 344866 309966 344898
rect 311378 345454 311618 345486
rect 311378 345218 311380 345454
rect 311616 345218 311618 345454
rect 311378 345134 311618 345218
rect 311378 344898 311380 345134
rect 311616 344898 311618 345134
rect 311378 344866 311618 344898
rect 312184 345454 312424 345486
rect 312184 345218 312186 345454
rect 312422 345218 312424 345454
rect 312184 345134 312424 345218
rect 312184 344898 312186 345134
rect 312422 344898 312424 345134
rect 312184 344866 312424 344898
rect 321184 345454 321424 345486
rect 321184 345218 321186 345454
rect 321422 345218 321424 345454
rect 321184 345134 321424 345218
rect 321184 344898 321186 345134
rect 321422 344898 321424 345134
rect 321184 344866 321424 344898
rect 330184 345454 330424 345486
rect 330184 345218 330186 345454
rect 330422 345218 330424 345454
rect 330184 345134 330424 345218
rect 330184 344898 330186 345134
rect 330422 344898 330424 345134
rect 330184 344866 330424 344898
rect 339184 345454 339424 345486
rect 339184 345218 339186 345454
rect 339422 345218 339424 345454
rect 339184 345134 339424 345218
rect 339184 344898 339186 345134
rect 339422 344898 339424 345134
rect 339184 344866 339424 344898
rect 348184 345454 348424 345486
rect 348184 345218 348186 345454
rect 348422 345218 348424 345454
rect 348184 345134 348424 345218
rect 348184 344898 348186 345134
rect 348422 344898 348424 345134
rect 348184 344866 348424 344898
rect 350746 345454 350986 345486
rect 350746 345218 350748 345454
rect 350984 345218 350986 345454
rect 350746 345134 350986 345218
rect 350746 344898 350748 345134
rect 350984 344898 350986 345134
rect 350746 344866 350986 344898
rect 352398 345454 352638 345486
rect 352398 345218 352400 345454
rect 352636 345218 352638 345454
rect 352398 345134 352638 345218
rect 352398 344898 352400 345134
rect 352636 344898 352638 345134
rect 352398 344866 352638 344898
rect 353204 345454 353444 345486
rect 353204 345218 353206 345454
rect 353442 345218 353444 345454
rect 353204 345134 353444 345218
rect 353204 344898 353206 345134
rect 353442 344898 353444 345134
rect 353204 344866 353444 344898
rect 362204 345454 362444 345486
rect 362204 345218 362206 345454
rect 362442 345218 362444 345454
rect 362204 345134 362444 345218
rect 362204 344898 362206 345134
rect 362442 344898 362444 345134
rect 362204 344866 362444 344898
rect 371204 345454 371444 345486
rect 371204 345218 371206 345454
rect 371442 345218 371444 345454
rect 371204 345134 371444 345218
rect 371204 344898 371206 345134
rect 371442 344898 371444 345134
rect 371204 344866 371444 344898
rect 380204 345454 380444 345486
rect 380204 345218 380206 345454
rect 380442 345218 380444 345454
rect 380204 345134 380444 345218
rect 380204 344898 380206 345134
rect 380442 344898 380444 345134
rect 380204 344866 380444 344898
rect 389204 345454 389444 345486
rect 389204 345218 389206 345454
rect 389442 345218 389444 345454
rect 389204 345134 389444 345218
rect 389204 344898 389206 345134
rect 389442 344898 389444 345134
rect 389204 344866 389444 344898
rect 391766 345454 392006 345486
rect 391766 345218 391768 345454
rect 392004 345218 392006 345454
rect 391766 345134 392006 345218
rect 391766 344898 391768 345134
rect 392004 344898 392006 345134
rect 391766 344866 392006 344898
rect 392418 345454 392658 345486
rect 392418 345218 392420 345454
rect 392656 345218 392658 345454
rect 392418 345134 392658 345218
rect 392418 344898 392420 345134
rect 392656 344898 392658 345134
rect 392418 344866 392658 344898
rect 393224 345454 393464 345486
rect 393224 345218 393226 345454
rect 393462 345218 393464 345454
rect 393224 345134 393464 345218
rect 393224 344898 393226 345134
rect 393462 344898 393464 345134
rect 393224 344866 393464 344898
rect 402224 345454 402464 345486
rect 402224 345218 402226 345454
rect 402462 345218 402464 345454
rect 402224 345134 402464 345218
rect 402224 344898 402226 345134
rect 402462 344898 402464 345134
rect 402224 344866 402464 344898
rect 411224 345454 411464 345486
rect 411224 345218 411226 345454
rect 411462 345218 411464 345454
rect 411224 345134 411464 345218
rect 411224 344898 411226 345134
rect 411462 344898 411464 345134
rect 411224 344866 411464 344898
rect 420224 345454 420464 345486
rect 420224 345218 420226 345454
rect 420462 345218 420464 345454
rect 420224 345134 420464 345218
rect 420224 344898 420226 345134
rect 420462 344898 420464 345134
rect 420224 344866 420464 344898
rect 429224 345454 429464 345486
rect 429224 345218 429226 345454
rect 429462 345218 429464 345454
rect 429224 345134 429464 345218
rect 429224 344898 429226 345134
rect 429462 344898 429464 345134
rect 429224 344866 429464 344898
rect 431786 345454 432026 345486
rect 431786 345218 431788 345454
rect 432024 345218 432026 345454
rect 431786 345134 432026 345218
rect 431786 344898 431788 345134
rect 432024 344898 432026 345134
rect 431786 344866 432026 344898
rect 432438 345454 432678 345486
rect 432438 345218 432440 345454
rect 432676 345218 432678 345454
rect 432438 345134 432678 345218
rect 432438 344898 432440 345134
rect 432676 344898 432678 345134
rect 432438 344866 432678 344898
rect 433244 345454 433484 345486
rect 433244 345218 433246 345454
rect 433482 345218 433484 345454
rect 433244 345134 433484 345218
rect 433244 344898 433246 345134
rect 433482 344898 433484 345134
rect 433244 344866 433484 344898
rect 439790 345454 440030 345486
rect 439790 345218 439792 345454
rect 440028 345218 440030 345454
rect 439790 345134 440030 345218
rect 439790 344898 439792 345134
rect 440028 344898 440030 345134
rect 439790 344866 440030 344898
rect 457008 345454 457248 345486
rect 457008 345218 457010 345454
rect 457246 345218 457248 345454
rect 457008 345134 457248 345218
rect 457008 344898 457010 345134
rect 457246 344898 457248 345134
rect 457008 344866 457248 344898
rect 579288 345454 579888 345486
rect 579288 345218 579470 345454
rect 579706 345218 579888 345454
rect 579288 345134 579888 345218
rect 579288 344898 579470 345134
rect 579706 344898 579888 345134
rect 579288 344866 579888 344898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect 5200 327454 5800 327486
rect 5200 327218 5382 327454
rect 5618 327218 5800 327454
rect 5200 327134 5800 327218
rect 5200 326898 5382 327134
rect 5618 326898 5800 327134
rect 5200 326866 5800 326898
rect 127456 327454 127696 327486
rect 127456 327218 127458 327454
rect 127694 327218 127696 327454
rect 127456 327134 127696 327218
rect 127456 326898 127458 327134
rect 127694 326898 127696 327134
rect 127456 326866 127696 326898
rect 140654 327454 140894 327486
rect 140654 327218 140656 327454
rect 140892 327218 140894 327454
rect 140654 327134 140894 327218
rect 140654 326898 140656 327134
rect 140892 326898 140894 327134
rect 140654 326866 140894 326898
rect 141500 327454 141740 327486
rect 141500 327218 141502 327454
rect 141738 327218 141740 327454
rect 141500 327134 141740 327218
rect 141500 326898 141502 327134
rect 141738 326898 141740 327134
rect 141500 326866 141740 326898
rect 147286 327454 147526 327486
rect 147286 327218 147288 327454
rect 147524 327218 147526 327454
rect 147286 327134 147526 327218
rect 147286 326898 147288 327134
rect 147524 326898 147526 327134
rect 147286 326866 147526 326898
rect 149658 327454 149898 327486
rect 149658 327218 149660 327454
rect 149896 327218 149898 327454
rect 149658 327134 149898 327218
rect 149658 326898 149660 327134
rect 149896 326898 149898 327134
rect 149658 326866 149898 326898
rect 150504 327454 150744 327486
rect 150504 327218 150506 327454
rect 150742 327218 150744 327454
rect 150504 327134 150744 327218
rect 150504 326898 150506 327134
rect 150742 326898 150744 327134
rect 150504 326866 150744 326898
rect 159504 327454 159744 327486
rect 159504 327218 159506 327454
rect 159742 327218 159744 327454
rect 159504 327134 159744 327218
rect 159504 326898 159506 327134
rect 159742 326898 159744 327134
rect 159504 326866 159744 326898
rect 168504 327454 168744 327486
rect 168504 327218 168506 327454
rect 168742 327218 168744 327454
rect 168504 327134 168744 327218
rect 168504 326898 168506 327134
rect 168742 326898 168744 327134
rect 168504 326866 168744 326898
rect 177504 327454 177744 327486
rect 177504 327218 177506 327454
rect 177742 327218 177744 327454
rect 177504 327134 177744 327218
rect 177504 326898 177506 327134
rect 177742 326898 177744 327134
rect 177504 326866 177744 326898
rect 186504 327454 186744 327486
rect 186504 327218 186506 327454
rect 186742 327218 186744 327454
rect 186504 327134 186744 327218
rect 186504 326898 186506 327134
rect 186742 326898 186744 327134
rect 186504 326866 186744 326898
rect 188306 327454 188546 327486
rect 188306 327218 188308 327454
rect 188544 327218 188546 327454
rect 188306 327134 188546 327218
rect 188306 326898 188308 327134
rect 188544 326898 188546 327134
rect 188306 326866 188546 326898
rect 189766 327454 190006 327486
rect 189766 327218 189768 327454
rect 190004 327218 190006 327454
rect 189766 327134 190006 327218
rect 189766 326898 189768 327134
rect 190004 326898 190006 327134
rect 189766 326866 190006 326898
rect 190678 327454 190918 327486
rect 190678 327218 190680 327454
rect 190916 327218 190918 327454
rect 190678 327134 190918 327218
rect 190678 326898 190680 327134
rect 190916 326898 190918 327134
rect 190678 326866 190918 326898
rect 191524 327454 191764 327486
rect 191524 327218 191526 327454
rect 191762 327218 191764 327454
rect 191524 327134 191764 327218
rect 191524 326898 191526 327134
rect 191762 326898 191764 327134
rect 191524 326866 191764 326898
rect 200524 327454 200764 327486
rect 200524 327218 200526 327454
rect 200762 327218 200764 327454
rect 200524 327134 200764 327218
rect 200524 326898 200526 327134
rect 200762 326898 200764 327134
rect 200524 326866 200764 326898
rect 209524 327454 209764 327486
rect 209524 327218 209526 327454
rect 209762 327218 209764 327454
rect 209524 327134 209764 327218
rect 209524 326898 209526 327134
rect 209762 326898 209764 327134
rect 209524 326866 209764 326898
rect 218524 327454 218764 327486
rect 218524 327218 218526 327454
rect 218762 327218 218764 327454
rect 218524 327134 218764 327218
rect 218524 326898 218526 327134
rect 218762 326898 218764 327134
rect 218524 326866 218764 326898
rect 227524 327454 227764 327486
rect 227524 327218 227526 327454
rect 227762 327218 227764 327454
rect 227524 327134 227764 327218
rect 227524 326898 227526 327134
rect 227762 326898 227764 327134
rect 227524 326866 227764 326898
rect 229326 327454 229566 327486
rect 229326 327218 229328 327454
rect 229564 327218 229566 327454
rect 229326 327134 229566 327218
rect 229326 326898 229328 327134
rect 229564 326898 229566 327134
rect 229326 326866 229566 326898
rect 230698 327454 230938 327486
rect 230698 327218 230700 327454
rect 230936 327218 230938 327454
rect 230698 327134 230938 327218
rect 230698 326898 230700 327134
rect 230936 326898 230938 327134
rect 230698 326866 230938 326898
rect 231544 327454 231784 327486
rect 231544 327218 231546 327454
rect 231782 327218 231784 327454
rect 231544 327134 231784 327218
rect 231544 326898 231546 327134
rect 231782 326898 231784 327134
rect 231544 326866 231784 326898
rect 240544 327454 240784 327486
rect 240544 327218 240546 327454
rect 240782 327218 240784 327454
rect 240544 327134 240784 327218
rect 240544 326898 240546 327134
rect 240782 326898 240784 327134
rect 240544 326866 240784 326898
rect 249544 327454 249784 327486
rect 249544 327218 249546 327454
rect 249782 327218 249784 327454
rect 249544 327134 249784 327218
rect 249544 326898 249546 327134
rect 249782 326898 249784 327134
rect 249544 326866 249784 326898
rect 258544 327454 258784 327486
rect 258544 327218 258546 327454
rect 258782 327218 258784 327454
rect 258544 327134 258784 327218
rect 258544 326898 258546 327134
rect 258782 326898 258784 327134
rect 258544 326866 258784 326898
rect 267544 327454 267784 327486
rect 267544 327218 267546 327454
rect 267782 327218 267784 327454
rect 267544 327134 267784 327218
rect 267544 326898 267546 327134
rect 267782 326898 267784 327134
rect 267544 326866 267784 326898
rect 269346 327454 269586 327486
rect 269346 327218 269348 327454
rect 269584 327218 269586 327454
rect 269346 327134 269586 327218
rect 269346 326898 269348 327134
rect 269584 326898 269586 327134
rect 269346 326866 269586 326898
rect 270718 327454 270958 327486
rect 270718 327218 270720 327454
rect 270956 327218 270958 327454
rect 270718 327134 270958 327218
rect 270718 326898 270720 327134
rect 270956 326898 270958 327134
rect 270718 326866 270958 326898
rect 271564 327454 271804 327486
rect 271564 327218 271566 327454
rect 271802 327218 271804 327454
rect 271564 327134 271804 327218
rect 271564 326898 271566 327134
rect 271802 326898 271804 327134
rect 271564 326866 271804 326898
rect 280564 327454 280804 327486
rect 280564 327218 280566 327454
rect 280802 327218 280804 327454
rect 280564 327134 280804 327218
rect 280564 326898 280566 327134
rect 280802 326898 280804 327134
rect 280564 326866 280804 326898
rect 289564 327454 289804 327486
rect 289564 327218 289566 327454
rect 289802 327218 289804 327454
rect 289564 327134 289804 327218
rect 289564 326898 289566 327134
rect 289802 326898 289804 327134
rect 289564 326866 289804 326898
rect 298564 327454 298804 327486
rect 298564 327218 298566 327454
rect 298802 327218 298804 327454
rect 298564 327134 298804 327218
rect 298564 326898 298566 327134
rect 298802 326898 298804 327134
rect 298564 326866 298804 326898
rect 307564 327454 307804 327486
rect 307564 327218 307566 327454
rect 307802 327218 307804 327454
rect 307564 327134 307804 327218
rect 307564 326898 307566 327134
rect 307802 326898 307804 327134
rect 307564 326866 307804 326898
rect 309366 327454 309606 327486
rect 309366 327218 309368 327454
rect 309604 327218 309606 327454
rect 309366 327134 309606 327218
rect 309366 326898 309368 327134
rect 309604 326898 309606 327134
rect 309366 326866 309606 326898
rect 311738 327454 311978 327486
rect 311738 327218 311740 327454
rect 311976 327218 311978 327454
rect 311738 327134 311978 327218
rect 311738 326898 311740 327134
rect 311976 326898 311978 327134
rect 311738 326866 311978 326898
rect 312584 327454 312824 327486
rect 312584 327218 312586 327454
rect 312822 327218 312824 327454
rect 312584 327134 312824 327218
rect 312584 326898 312586 327134
rect 312822 326898 312824 327134
rect 312584 326866 312824 326898
rect 321584 327454 321824 327486
rect 321584 327218 321586 327454
rect 321822 327218 321824 327454
rect 321584 327134 321824 327218
rect 321584 326898 321586 327134
rect 321822 326898 321824 327134
rect 321584 326866 321824 326898
rect 330584 327454 330824 327486
rect 330584 327218 330586 327454
rect 330822 327218 330824 327454
rect 330584 327134 330824 327218
rect 330584 326898 330586 327134
rect 330822 326898 330824 327134
rect 330584 326866 330824 326898
rect 339584 327454 339824 327486
rect 339584 327218 339586 327454
rect 339822 327218 339824 327454
rect 339584 327134 339824 327218
rect 339584 326898 339586 327134
rect 339822 326898 339824 327134
rect 339584 326866 339824 326898
rect 348584 327454 348824 327486
rect 348584 327218 348586 327454
rect 348822 327218 348824 327454
rect 348584 327134 348824 327218
rect 348584 326898 348586 327134
rect 348822 326898 348824 327134
rect 348584 326866 348824 326898
rect 350386 327454 350626 327486
rect 350386 327218 350388 327454
rect 350624 327218 350626 327454
rect 350386 327134 350626 327218
rect 350386 326898 350388 327134
rect 350624 326898 350626 327134
rect 350386 326866 350626 326898
rect 352758 327454 352998 327486
rect 352758 327218 352760 327454
rect 352996 327218 352998 327454
rect 352758 327134 352998 327218
rect 352758 326898 352760 327134
rect 352996 326898 352998 327134
rect 352758 326866 352998 326898
rect 353604 327454 353844 327486
rect 353604 327218 353606 327454
rect 353842 327218 353844 327454
rect 353604 327134 353844 327218
rect 353604 326898 353606 327134
rect 353842 326898 353844 327134
rect 353604 326866 353844 326898
rect 362604 327454 362844 327486
rect 362604 327218 362606 327454
rect 362842 327218 362844 327454
rect 362604 327134 362844 327218
rect 362604 326898 362606 327134
rect 362842 326898 362844 327134
rect 362604 326866 362844 326898
rect 371604 327454 371844 327486
rect 371604 327218 371606 327454
rect 371842 327218 371844 327454
rect 371604 327134 371844 327218
rect 371604 326898 371606 327134
rect 371842 326898 371844 327134
rect 371604 326866 371844 326898
rect 380604 327454 380844 327486
rect 380604 327218 380606 327454
rect 380842 327218 380844 327454
rect 380604 327134 380844 327218
rect 380604 326898 380606 327134
rect 380842 326898 380844 327134
rect 380604 326866 380844 326898
rect 389604 327454 389844 327486
rect 389604 327218 389606 327454
rect 389842 327218 389844 327454
rect 389604 327134 389844 327218
rect 389604 326898 389606 327134
rect 389842 326898 389844 327134
rect 389604 326866 389844 326898
rect 391406 327454 391646 327486
rect 391406 327218 391408 327454
rect 391644 327218 391646 327454
rect 391406 327134 391646 327218
rect 391406 326898 391408 327134
rect 391644 326898 391646 327134
rect 391406 326866 391646 326898
rect 392778 327454 393018 327486
rect 392778 327218 392780 327454
rect 393016 327218 393018 327454
rect 392778 327134 393018 327218
rect 392778 326898 392780 327134
rect 393016 326898 393018 327134
rect 392778 326866 393018 326898
rect 393624 327454 393864 327486
rect 393624 327218 393626 327454
rect 393862 327218 393864 327454
rect 393624 327134 393864 327218
rect 393624 326898 393626 327134
rect 393862 326898 393864 327134
rect 393624 326866 393864 326898
rect 402624 327454 402864 327486
rect 402624 327218 402626 327454
rect 402862 327218 402864 327454
rect 402624 327134 402864 327218
rect 402624 326898 402626 327134
rect 402862 326898 402864 327134
rect 402624 326866 402864 326898
rect 411624 327454 411864 327486
rect 411624 327218 411626 327454
rect 411862 327218 411864 327454
rect 411624 327134 411864 327218
rect 411624 326898 411626 327134
rect 411862 326898 411864 327134
rect 411624 326866 411864 326898
rect 420624 327454 420864 327486
rect 420624 327218 420626 327454
rect 420862 327218 420864 327454
rect 420624 327134 420864 327218
rect 420624 326898 420626 327134
rect 420862 326898 420864 327134
rect 420624 326866 420864 326898
rect 429624 327454 429864 327486
rect 429624 327218 429626 327454
rect 429862 327218 429864 327454
rect 429624 327134 429864 327218
rect 429624 326898 429626 327134
rect 429862 326898 429864 327134
rect 429624 326866 429864 326898
rect 431426 327454 431666 327486
rect 431426 327218 431428 327454
rect 431664 327218 431666 327454
rect 431426 327134 431666 327218
rect 431426 326898 431428 327134
rect 431664 326898 431666 327134
rect 431426 326866 431666 326898
rect 432798 327454 433038 327486
rect 432798 327218 432800 327454
rect 433036 327218 433038 327454
rect 432798 327134 433038 327218
rect 432798 326898 432800 327134
rect 433036 326898 433038 327134
rect 432798 326866 433038 326898
rect 433644 327454 433884 327486
rect 433644 327218 433646 327454
rect 433882 327218 433884 327454
rect 433644 327134 433884 327218
rect 433644 326898 433646 327134
rect 433882 326898 433884 327134
rect 433644 326866 433884 326898
rect 439430 327454 439670 327486
rect 439430 327218 439432 327454
rect 439668 327218 439670 327454
rect 439430 327134 439670 327218
rect 439430 326898 439432 327134
rect 439668 326898 439670 327134
rect 439430 326866 439670 326898
rect 456608 327454 456848 327486
rect 456608 327218 456610 327454
rect 456846 327218 456848 327454
rect 456608 327134 456848 327218
rect 456608 326898 456610 327134
rect 456846 326898 456848 327134
rect 456608 326866 456848 326898
rect 578488 327454 579088 327486
rect 578488 327218 578670 327454
rect 578906 327218 579088 327454
rect 578488 327134 579088 327218
rect 578488 326898 578670 327134
rect 578906 326898 579088 327134
rect 578488 326866 579088 326898
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 4400 309454 5000 309486
rect 4400 309218 4582 309454
rect 4818 309218 5000 309454
rect 4400 309134 5000 309218
rect 4400 308898 4582 309134
rect 4818 308898 5000 309134
rect 4400 308866 5000 308898
rect 127056 309454 127296 309486
rect 127056 309218 127058 309454
rect 127294 309218 127296 309454
rect 127056 309134 127296 309218
rect 127056 308898 127058 309134
rect 127294 308898 127296 309134
rect 127056 308866 127296 308898
rect 140294 309454 140534 309486
rect 140294 309218 140296 309454
rect 140532 309218 140534 309454
rect 140294 309134 140534 309218
rect 140294 308898 140296 309134
rect 140532 308898 140534 309134
rect 140294 308866 140534 308898
rect 141100 309454 141340 309486
rect 141100 309218 141102 309454
rect 141338 309218 141340 309454
rect 141100 309134 141340 309218
rect 141100 308898 141102 309134
rect 141338 308898 141340 309134
rect 141100 308866 141340 308898
rect 147646 309454 147886 309486
rect 147646 309218 147648 309454
rect 147884 309218 147886 309454
rect 147646 309134 147886 309218
rect 147646 308898 147648 309134
rect 147884 308898 147886 309134
rect 147646 308866 147886 308898
rect 149298 309454 149538 309486
rect 149298 309218 149300 309454
rect 149536 309218 149538 309454
rect 149298 309134 149538 309218
rect 149298 308898 149300 309134
rect 149536 308898 149538 309134
rect 149298 308866 149538 308898
rect 150104 309454 150344 309486
rect 150104 309218 150106 309454
rect 150342 309218 150344 309454
rect 150104 309134 150344 309218
rect 150104 308898 150106 309134
rect 150342 308898 150344 309134
rect 150104 308866 150344 308898
rect 159104 309454 159344 309486
rect 159104 309218 159106 309454
rect 159342 309218 159344 309454
rect 159104 309134 159344 309218
rect 159104 308898 159106 309134
rect 159342 308898 159344 309134
rect 159104 308866 159344 308898
rect 168104 309454 168344 309486
rect 168104 309218 168106 309454
rect 168342 309218 168344 309454
rect 168104 309134 168344 309218
rect 168104 308898 168106 309134
rect 168342 308898 168344 309134
rect 168104 308866 168344 308898
rect 177104 309454 177344 309486
rect 177104 309218 177106 309454
rect 177342 309218 177344 309454
rect 177104 309134 177344 309218
rect 177104 308898 177106 309134
rect 177342 308898 177344 309134
rect 177104 308866 177344 308898
rect 186104 309454 186344 309486
rect 186104 309218 186106 309454
rect 186342 309218 186344 309454
rect 186104 309134 186344 309218
rect 186104 308898 186106 309134
rect 186342 308898 186344 309134
rect 186104 308866 186344 308898
rect 188666 309454 188906 309486
rect 188666 309218 188668 309454
rect 188904 309218 188906 309454
rect 188666 309134 188906 309218
rect 188666 308898 188668 309134
rect 188904 308898 188906 309134
rect 188666 308866 188906 308898
rect 190318 309454 190558 309486
rect 190318 309218 190320 309454
rect 190556 309218 190558 309454
rect 190318 309134 190558 309218
rect 190318 308898 190320 309134
rect 190556 308898 190558 309134
rect 190318 308866 190558 308898
rect 191124 309454 191364 309486
rect 191124 309218 191126 309454
rect 191362 309218 191364 309454
rect 191124 309134 191364 309218
rect 191124 308898 191126 309134
rect 191362 308898 191364 309134
rect 191124 308866 191364 308898
rect 200124 309454 200364 309486
rect 200124 309218 200126 309454
rect 200362 309218 200364 309454
rect 200124 309134 200364 309218
rect 200124 308898 200126 309134
rect 200362 308898 200364 309134
rect 200124 308866 200364 308898
rect 209124 309454 209364 309486
rect 209124 309218 209126 309454
rect 209362 309218 209364 309454
rect 209124 309134 209364 309218
rect 209124 308898 209126 309134
rect 209362 308898 209364 309134
rect 209124 308866 209364 308898
rect 218124 309454 218364 309486
rect 218124 309218 218126 309454
rect 218362 309218 218364 309454
rect 218124 309134 218364 309218
rect 218124 308898 218126 309134
rect 218362 308898 218364 309134
rect 218124 308866 218364 308898
rect 227124 309454 227364 309486
rect 227124 309218 227126 309454
rect 227362 309218 227364 309454
rect 227124 309134 227364 309218
rect 227124 308898 227126 309134
rect 227362 308898 227364 309134
rect 227124 308866 227364 308898
rect 229686 309454 229926 309486
rect 229686 309218 229688 309454
rect 229924 309218 229926 309454
rect 229686 309134 229926 309218
rect 229686 308898 229688 309134
rect 229924 308898 229926 309134
rect 229686 308866 229926 308898
rect 230338 309454 230578 309486
rect 230338 309218 230340 309454
rect 230576 309218 230578 309454
rect 230338 309134 230578 309218
rect 230338 308898 230340 309134
rect 230576 308898 230578 309134
rect 230338 308866 230578 308898
rect 231144 309454 231384 309486
rect 231144 309218 231146 309454
rect 231382 309218 231384 309454
rect 231144 309134 231384 309218
rect 231144 308898 231146 309134
rect 231382 308898 231384 309134
rect 231144 308866 231384 308898
rect 240144 309454 240384 309486
rect 240144 309218 240146 309454
rect 240382 309218 240384 309454
rect 240144 309134 240384 309218
rect 240144 308898 240146 309134
rect 240382 308898 240384 309134
rect 240144 308866 240384 308898
rect 249144 309454 249384 309486
rect 249144 309218 249146 309454
rect 249382 309218 249384 309454
rect 249144 309134 249384 309218
rect 249144 308898 249146 309134
rect 249382 308898 249384 309134
rect 249144 308866 249384 308898
rect 258144 309454 258384 309486
rect 258144 309218 258146 309454
rect 258382 309218 258384 309454
rect 258144 309134 258384 309218
rect 258144 308898 258146 309134
rect 258382 308898 258384 309134
rect 258144 308866 258384 308898
rect 267144 309454 267384 309486
rect 267144 309218 267146 309454
rect 267382 309218 267384 309454
rect 267144 309134 267384 309218
rect 267144 308898 267146 309134
rect 267382 308898 267384 309134
rect 267144 308866 267384 308898
rect 269706 309454 269946 309486
rect 269706 309218 269708 309454
rect 269944 309218 269946 309454
rect 269706 309134 269946 309218
rect 269706 308898 269708 309134
rect 269944 308898 269946 309134
rect 269706 308866 269946 308898
rect 270358 309454 270598 309486
rect 270358 309218 270360 309454
rect 270596 309218 270598 309454
rect 270358 309134 270598 309218
rect 270358 308898 270360 309134
rect 270596 308898 270598 309134
rect 270358 308866 270598 308898
rect 271164 309454 271404 309486
rect 271164 309218 271166 309454
rect 271402 309218 271404 309454
rect 271164 309134 271404 309218
rect 271164 308898 271166 309134
rect 271402 308898 271404 309134
rect 271164 308866 271404 308898
rect 280164 309454 280404 309486
rect 280164 309218 280166 309454
rect 280402 309218 280404 309454
rect 280164 309134 280404 309218
rect 280164 308898 280166 309134
rect 280402 308898 280404 309134
rect 280164 308866 280404 308898
rect 289164 309454 289404 309486
rect 289164 309218 289166 309454
rect 289402 309218 289404 309454
rect 289164 309134 289404 309218
rect 289164 308898 289166 309134
rect 289402 308898 289404 309134
rect 289164 308866 289404 308898
rect 298164 309454 298404 309486
rect 298164 309218 298166 309454
rect 298402 309218 298404 309454
rect 298164 309134 298404 309218
rect 298164 308898 298166 309134
rect 298402 308898 298404 309134
rect 298164 308866 298404 308898
rect 307164 309454 307404 309486
rect 307164 309218 307166 309454
rect 307402 309218 307404 309454
rect 307164 309134 307404 309218
rect 307164 308898 307166 309134
rect 307402 308898 307404 309134
rect 307164 308866 307404 308898
rect 309726 309454 309966 309486
rect 309726 309218 309728 309454
rect 309964 309218 309966 309454
rect 309726 309134 309966 309218
rect 309726 308898 309728 309134
rect 309964 308898 309966 309134
rect 309726 308866 309966 308898
rect 311378 309454 311618 309486
rect 311378 309218 311380 309454
rect 311616 309218 311618 309454
rect 311378 309134 311618 309218
rect 311378 308898 311380 309134
rect 311616 308898 311618 309134
rect 311378 308866 311618 308898
rect 312184 309454 312424 309486
rect 312184 309218 312186 309454
rect 312422 309218 312424 309454
rect 312184 309134 312424 309218
rect 312184 308898 312186 309134
rect 312422 308898 312424 309134
rect 312184 308866 312424 308898
rect 321184 309454 321424 309486
rect 321184 309218 321186 309454
rect 321422 309218 321424 309454
rect 321184 309134 321424 309218
rect 321184 308898 321186 309134
rect 321422 308898 321424 309134
rect 321184 308866 321424 308898
rect 330184 309454 330424 309486
rect 330184 309218 330186 309454
rect 330422 309218 330424 309454
rect 330184 309134 330424 309218
rect 330184 308898 330186 309134
rect 330422 308898 330424 309134
rect 330184 308866 330424 308898
rect 339184 309454 339424 309486
rect 339184 309218 339186 309454
rect 339422 309218 339424 309454
rect 339184 309134 339424 309218
rect 339184 308898 339186 309134
rect 339422 308898 339424 309134
rect 339184 308866 339424 308898
rect 348184 309454 348424 309486
rect 348184 309218 348186 309454
rect 348422 309218 348424 309454
rect 348184 309134 348424 309218
rect 348184 308898 348186 309134
rect 348422 308898 348424 309134
rect 348184 308866 348424 308898
rect 350746 309454 350986 309486
rect 350746 309218 350748 309454
rect 350984 309218 350986 309454
rect 350746 309134 350986 309218
rect 350746 308898 350748 309134
rect 350984 308898 350986 309134
rect 350746 308866 350986 308898
rect 352398 309454 352638 309486
rect 352398 309218 352400 309454
rect 352636 309218 352638 309454
rect 352398 309134 352638 309218
rect 352398 308898 352400 309134
rect 352636 308898 352638 309134
rect 352398 308866 352638 308898
rect 353204 309454 353444 309486
rect 353204 309218 353206 309454
rect 353442 309218 353444 309454
rect 353204 309134 353444 309218
rect 353204 308898 353206 309134
rect 353442 308898 353444 309134
rect 353204 308866 353444 308898
rect 362204 309454 362444 309486
rect 362204 309218 362206 309454
rect 362442 309218 362444 309454
rect 362204 309134 362444 309218
rect 362204 308898 362206 309134
rect 362442 308898 362444 309134
rect 362204 308866 362444 308898
rect 371204 309454 371444 309486
rect 371204 309218 371206 309454
rect 371442 309218 371444 309454
rect 371204 309134 371444 309218
rect 371204 308898 371206 309134
rect 371442 308898 371444 309134
rect 371204 308866 371444 308898
rect 380204 309454 380444 309486
rect 380204 309218 380206 309454
rect 380442 309218 380444 309454
rect 380204 309134 380444 309218
rect 380204 308898 380206 309134
rect 380442 308898 380444 309134
rect 380204 308866 380444 308898
rect 389204 309454 389444 309486
rect 389204 309218 389206 309454
rect 389442 309218 389444 309454
rect 389204 309134 389444 309218
rect 389204 308898 389206 309134
rect 389442 308898 389444 309134
rect 389204 308866 389444 308898
rect 391766 309454 392006 309486
rect 391766 309218 391768 309454
rect 392004 309218 392006 309454
rect 391766 309134 392006 309218
rect 391766 308898 391768 309134
rect 392004 308898 392006 309134
rect 391766 308866 392006 308898
rect 392418 309454 392658 309486
rect 392418 309218 392420 309454
rect 392656 309218 392658 309454
rect 392418 309134 392658 309218
rect 392418 308898 392420 309134
rect 392656 308898 392658 309134
rect 392418 308866 392658 308898
rect 393224 309454 393464 309486
rect 393224 309218 393226 309454
rect 393462 309218 393464 309454
rect 393224 309134 393464 309218
rect 393224 308898 393226 309134
rect 393462 308898 393464 309134
rect 393224 308866 393464 308898
rect 402224 309454 402464 309486
rect 402224 309218 402226 309454
rect 402462 309218 402464 309454
rect 402224 309134 402464 309218
rect 402224 308898 402226 309134
rect 402462 308898 402464 309134
rect 402224 308866 402464 308898
rect 411224 309454 411464 309486
rect 411224 309218 411226 309454
rect 411462 309218 411464 309454
rect 411224 309134 411464 309218
rect 411224 308898 411226 309134
rect 411462 308898 411464 309134
rect 411224 308866 411464 308898
rect 420224 309454 420464 309486
rect 420224 309218 420226 309454
rect 420462 309218 420464 309454
rect 420224 309134 420464 309218
rect 420224 308898 420226 309134
rect 420462 308898 420464 309134
rect 420224 308866 420464 308898
rect 429224 309454 429464 309486
rect 429224 309218 429226 309454
rect 429462 309218 429464 309454
rect 429224 309134 429464 309218
rect 429224 308898 429226 309134
rect 429462 308898 429464 309134
rect 429224 308866 429464 308898
rect 431786 309454 432026 309486
rect 431786 309218 431788 309454
rect 432024 309218 432026 309454
rect 431786 309134 432026 309218
rect 431786 308898 431788 309134
rect 432024 308898 432026 309134
rect 431786 308866 432026 308898
rect 432438 309454 432678 309486
rect 432438 309218 432440 309454
rect 432676 309218 432678 309454
rect 432438 309134 432678 309218
rect 432438 308898 432440 309134
rect 432676 308898 432678 309134
rect 432438 308866 432678 308898
rect 433244 309454 433484 309486
rect 433244 309218 433246 309454
rect 433482 309218 433484 309454
rect 433244 309134 433484 309218
rect 433244 308898 433246 309134
rect 433482 308898 433484 309134
rect 433244 308866 433484 308898
rect 439790 309454 440030 309486
rect 439790 309218 439792 309454
rect 440028 309218 440030 309454
rect 439790 309134 440030 309218
rect 439790 308898 439792 309134
rect 440028 308898 440030 309134
rect 439790 308866 440030 308898
rect 457008 309454 457248 309486
rect 457008 309218 457010 309454
rect 457246 309218 457248 309454
rect 457008 309134 457248 309218
rect 457008 308898 457010 309134
rect 457246 308898 457248 309134
rect 457008 308866 457248 308898
rect 579288 309454 579888 309486
rect 579288 309218 579470 309454
rect 579706 309218 579888 309454
rect 579288 309134 579888 309218
rect 579288 308898 579470 309134
rect 579706 308898 579888 309134
rect 579288 308866 579888 308898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect 5200 291454 5800 291486
rect 5200 291218 5382 291454
rect 5618 291218 5800 291454
rect 5200 291134 5800 291218
rect 5200 290898 5382 291134
rect 5618 290898 5800 291134
rect 5200 290866 5800 290898
rect 108638 291454 108878 291486
rect 108638 291218 108640 291454
rect 108876 291218 108878 291454
rect 108638 291134 108878 291218
rect 108638 290898 108640 291134
rect 108876 290898 108878 291134
rect 108638 290866 108878 290898
rect 109484 291454 109724 291486
rect 109484 291218 109486 291454
rect 109722 291218 109724 291454
rect 109484 291134 109724 291218
rect 109484 290898 109486 291134
rect 109722 290898 109724 291134
rect 109484 290866 109724 290898
rect 118484 291454 118724 291486
rect 118484 291218 118486 291454
rect 118722 291218 118724 291454
rect 118484 291134 118724 291218
rect 118484 290898 118486 291134
rect 118722 290898 118724 291134
rect 118484 290866 118724 290898
rect 127484 291454 127724 291486
rect 127484 291218 127486 291454
rect 127722 291218 127724 291454
rect 127484 291134 127724 291218
rect 127484 290898 127486 291134
rect 127722 290898 127724 291134
rect 127484 290866 127724 290898
rect 136484 291454 136724 291486
rect 136484 291218 136486 291454
rect 136722 291218 136724 291454
rect 136484 291134 136724 291218
rect 136484 290898 136486 291134
rect 136722 290898 136724 291134
rect 136484 290866 136724 290898
rect 145484 291454 145724 291486
rect 145484 291218 145486 291454
rect 145722 291218 145724 291454
rect 145484 291134 145724 291218
rect 145484 290898 145486 291134
rect 145722 290898 145724 291134
rect 145484 290866 145724 290898
rect 147286 291454 147526 291486
rect 147286 291218 147288 291454
rect 147524 291218 147526 291454
rect 147286 291134 147526 291218
rect 147286 290898 147288 291134
rect 147524 290898 147526 291134
rect 147286 290866 147526 290898
rect 149658 291454 149898 291486
rect 149658 291218 149660 291454
rect 149896 291218 149898 291454
rect 149658 291134 149898 291218
rect 149658 290898 149660 291134
rect 149896 290898 149898 291134
rect 149658 290866 149898 290898
rect 150504 291454 150744 291486
rect 150504 291218 150506 291454
rect 150742 291218 150744 291454
rect 150504 291134 150744 291218
rect 150504 290898 150506 291134
rect 150742 290898 150744 291134
rect 150504 290866 150744 290898
rect 159504 291454 159744 291486
rect 159504 291218 159506 291454
rect 159742 291218 159744 291454
rect 159504 291134 159744 291218
rect 159504 290898 159506 291134
rect 159742 290898 159744 291134
rect 159504 290866 159744 290898
rect 168504 291454 168744 291486
rect 168504 291218 168506 291454
rect 168742 291218 168744 291454
rect 168504 291134 168744 291218
rect 168504 290898 168506 291134
rect 168742 290898 168744 291134
rect 168504 290866 168744 290898
rect 177504 291454 177744 291486
rect 177504 291218 177506 291454
rect 177742 291218 177744 291454
rect 177504 291134 177744 291218
rect 177504 290898 177506 291134
rect 177742 290898 177744 291134
rect 177504 290866 177744 290898
rect 186504 291454 186744 291486
rect 186504 291218 186506 291454
rect 186742 291218 186744 291454
rect 186504 291134 186744 291218
rect 186504 290898 186506 291134
rect 186742 290898 186744 291134
rect 186504 290866 186744 290898
rect 188306 291454 188546 291486
rect 188306 291218 188308 291454
rect 188544 291218 188546 291454
rect 188306 291134 188546 291218
rect 188306 290898 188308 291134
rect 188544 290898 188546 291134
rect 188306 290866 188546 290898
rect 190678 291454 190918 291486
rect 190678 291218 190680 291454
rect 190916 291218 190918 291454
rect 190678 291134 190918 291218
rect 190678 290898 190680 291134
rect 190916 290898 190918 291134
rect 190678 290866 190918 290898
rect 191524 291454 191764 291486
rect 191524 291218 191526 291454
rect 191762 291218 191764 291454
rect 191524 291134 191764 291218
rect 191524 290898 191526 291134
rect 191762 290898 191764 291134
rect 191524 290866 191764 290898
rect 200524 291454 200764 291486
rect 200524 291218 200526 291454
rect 200762 291218 200764 291454
rect 200524 291134 200764 291218
rect 200524 290898 200526 291134
rect 200762 290898 200764 291134
rect 200524 290866 200764 290898
rect 209524 291454 209764 291486
rect 209524 291218 209526 291454
rect 209762 291218 209764 291454
rect 209524 291134 209764 291218
rect 209524 290898 209526 291134
rect 209762 290898 209764 291134
rect 209524 290866 209764 290898
rect 218524 291454 218764 291486
rect 218524 291218 218526 291454
rect 218762 291218 218764 291454
rect 218524 291134 218764 291218
rect 218524 290898 218526 291134
rect 218762 290898 218764 291134
rect 218524 290866 218764 290898
rect 227524 291454 227764 291486
rect 227524 291218 227526 291454
rect 227762 291218 227764 291454
rect 227524 291134 227764 291218
rect 227524 290898 227526 291134
rect 227762 290898 227764 291134
rect 227524 290866 227764 290898
rect 229326 291454 229566 291486
rect 229326 291218 229328 291454
rect 229564 291218 229566 291454
rect 229326 291134 229566 291218
rect 229326 290898 229328 291134
rect 229564 290898 229566 291134
rect 229326 290866 229566 290898
rect 230698 291454 230938 291486
rect 230698 291218 230700 291454
rect 230936 291218 230938 291454
rect 230698 291134 230938 291218
rect 230698 290898 230700 291134
rect 230936 290898 230938 291134
rect 230698 290866 230938 290898
rect 231544 291454 231784 291486
rect 231544 291218 231546 291454
rect 231782 291218 231784 291454
rect 231544 291134 231784 291218
rect 231544 290898 231546 291134
rect 231782 290898 231784 291134
rect 231544 290866 231784 290898
rect 240544 291454 240784 291486
rect 240544 291218 240546 291454
rect 240782 291218 240784 291454
rect 240544 291134 240784 291218
rect 240544 290898 240546 291134
rect 240782 290898 240784 291134
rect 240544 290866 240784 290898
rect 249544 291454 249784 291486
rect 249544 291218 249546 291454
rect 249782 291218 249784 291454
rect 249544 291134 249784 291218
rect 249544 290898 249546 291134
rect 249782 290898 249784 291134
rect 249544 290866 249784 290898
rect 258544 291454 258784 291486
rect 258544 291218 258546 291454
rect 258782 291218 258784 291454
rect 258544 291134 258784 291218
rect 258544 290898 258546 291134
rect 258782 290898 258784 291134
rect 258544 290866 258784 290898
rect 267544 291454 267784 291486
rect 267544 291218 267546 291454
rect 267782 291218 267784 291454
rect 267544 291134 267784 291218
rect 267544 290898 267546 291134
rect 267782 290898 267784 291134
rect 267544 290866 267784 290898
rect 269346 291454 269586 291486
rect 269346 291218 269348 291454
rect 269584 291218 269586 291454
rect 269346 291134 269586 291218
rect 269346 290898 269348 291134
rect 269584 290898 269586 291134
rect 269346 290866 269586 290898
rect 270718 291454 270958 291486
rect 270718 291218 270720 291454
rect 270956 291218 270958 291454
rect 270718 291134 270958 291218
rect 270718 290898 270720 291134
rect 270956 290898 270958 291134
rect 270718 290866 270958 290898
rect 271564 291454 271804 291486
rect 271564 291218 271566 291454
rect 271802 291218 271804 291454
rect 271564 291134 271804 291218
rect 271564 290898 271566 291134
rect 271802 290898 271804 291134
rect 271564 290866 271804 290898
rect 280564 291454 280804 291486
rect 280564 291218 280566 291454
rect 280802 291218 280804 291454
rect 280564 291134 280804 291218
rect 280564 290898 280566 291134
rect 280802 290898 280804 291134
rect 280564 290866 280804 290898
rect 289564 291454 289804 291486
rect 289564 291218 289566 291454
rect 289802 291218 289804 291454
rect 289564 291134 289804 291218
rect 289564 290898 289566 291134
rect 289802 290898 289804 291134
rect 289564 290866 289804 290898
rect 298564 291454 298804 291486
rect 298564 291218 298566 291454
rect 298802 291218 298804 291454
rect 298564 291134 298804 291218
rect 298564 290898 298566 291134
rect 298802 290898 298804 291134
rect 298564 290866 298804 290898
rect 307564 291454 307804 291486
rect 307564 291218 307566 291454
rect 307802 291218 307804 291454
rect 307564 291134 307804 291218
rect 307564 290898 307566 291134
rect 307802 290898 307804 291134
rect 307564 290866 307804 290898
rect 309366 291454 309606 291486
rect 309366 291218 309368 291454
rect 309604 291218 309606 291454
rect 309366 291134 309606 291218
rect 309366 290898 309368 291134
rect 309604 290898 309606 291134
rect 309366 290866 309606 290898
rect 311738 291454 311978 291486
rect 311738 291218 311740 291454
rect 311976 291218 311978 291454
rect 311738 291134 311978 291218
rect 311738 290898 311740 291134
rect 311976 290898 311978 291134
rect 311738 290866 311978 290898
rect 312584 291454 312824 291486
rect 312584 291218 312586 291454
rect 312822 291218 312824 291454
rect 312584 291134 312824 291218
rect 312584 290898 312586 291134
rect 312822 290898 312824 291134
rect 312584 290866 312824 290898
rect 321584 291454 321824 291486
rect 321584 291218 321586 291454
rect 321822 291218 321824 291454
rect 321584 291134 321824 291218
rect 321584 290898 321586 291134
rect 321822 290898 321824 291134
rect 321584 290866 321824 290898
rect 330584 291454 330824 291486
rect 330584 291218 330586 291454
rect 330822 291218 330824 291454
rect 330584 291134 330824 291218
rect 330584 290898 330586 291134
rect 330822 290898 330824 291134
rect 330584 290866 330824 290898
rect 339584 291454 339824 291486
rect 339584 291218 339586 291454
rect 339822 291218 339824 291454
rect 339584 291134 339824 291218
rect 339584 290898 339586 291134
rect 339822 290898 339824 291134
rect 339584 290866 339824 290898
rect 348584 291454 348824 291486
rect 348584 291218 348586 291454
rect 348822 291218 348824 291454
rect 348584 291134 348824 291218
rect 348584 290898 348586 291134
rect 348822 290898 348824 291134
rect 348584 290866 348824 290898
rect 350386 291454 350626 291486
rect 350386 291218 350388 291454
rect 350624 291218 350626 291454
rect 350386 291134 350626 291218
rect 350386 290898 350388 291134
rect 350624 290898 350626 291134
rect 350386 290866 350626 290898
rect 352758 291454 352998 291486
rect 352758 291218 352760 291454
rect 352996 291218 352998 291454
rect 352758 291134 352998 291218
rect 352758 290898 352760 291134
rect 352996 290898 352998 291134
rect 352758 290866 352998 290898
rect 353604 291454 353844 291486
rect 353604 291218 353606 291454
rect 353842 291218 353844 291454
rect 353604 291134 353844 291218
rect 353604 290898 353606 291134
rect 353842 290898 353844 291134
rect 353604 290866 353844 290898
rect 362604 291454 362844 291486
rect 362604 291218 362606 291454
rect 362842 291218 362844 291454
rect 362604 291134 362844 291218
rect 362604 290898 362606 291134
rect 362842 290898 362844 291134
rect 362604 290866 362844 290898
rect 371604 291454 371844 291486
rect 371604 291218 371606 291454
rect 371842 291218 371844 291454
rect 371604 291134 371844 291218
rect 371604 290898 371606 291134
rect 371842 290898 371844 291134
rect 371604 290866 371844 290898
rect 380604 291454 380844 291486
rect 380604 291218 380606 291454
rect 380842 291218 380844 291454
rect 380604 291134 380844 291218
rect 380604 290898 380606 291134
rect 380842 290898 380844 291134
rect 380604 290866 380844 290898
rect 389604 291454 389844 291486
rect 389604 291218 389606 291454
rect 389842 291218 389844 291454
rect 389604 291134 389844 291218
rect 389604 290898 389606 291134
rect 389842 290898 389844 291134
rect 389604 290866 389844 290898
rect 391406 291454 391646 291486
rect 391406 291218 391408 291454
rect 391644 291218 391646 291454
rect 391406 291134 391646 291218
rect 391406 290898 391408 291134
rect 391644 290898 391646 291134
rect 391406 290866 391646 290898
rect 392778 291454 393018 291486
rect 392778 291218 392780 291454
rect 393016 291218 393018 291454
rect 392778 291134 393018 291218
rect 392778 290898 392780 291134
rect 393016 290898 393018 291134
rect 392778 290866 393018 290898
rect 393624 291454 393864 291486
rect 393624 291218 393626 291454
rect 393862 291218 393864 291454
rect 393624 291134 393864 291218
rect 393624 290898 393626 291134
rect 393862 290898 393864 291134
rect 393624 290866 393864 290898
rect 402624 291454 402864 291486
rect 402624 291218 402626 291454
rect 402862 291218 402864 291454
rect 402624 291134 402864 291218
rect 402624 290898 402626 291134
rect 402862 290898 402864 291134
rect 402624 290866 402864 290898
rect 411624 291454 411864 291486
rect 411624 291218 411626 291454
rect 411862 291218 411864 291454
rect 411624 291134 411864 291218
rect 411624 290898 411626 291134
rect 411862 290898 411864 291134
rect 411624 290866 411864 290898
rect 420624 291454 420864 291486
rect 420624 291218 420626 291454
rect 420862 291218 420864 291454
rect 420624 291134 420864 291218
rect 420624 290898 420626 291134
rect 420862 290898 420864 291134
rect 420624 290866 420864 290898
rect 429624 291454 429864 291486
rect 429624 291218 429626 291454
rect 429862 291218 429864 291454
rect 429624 291134 429864 291218
rect 429624 290898 429626 291134
rect 429862 290898 429864 291134
rect 429624 290866 429864 290898
rect 431426 291454 431666 291486
rect 431426 291218 431428 291454
rect 431664 291218 431666 291454
rect 431426 291134 431666 291218
rect 431426 290898 431428 291134
rect 431664 290898 431666 291134
rect 431426 290866 431666 290898
rect 432798 291454 433038 291486
rect 432798 291218 432800 291454
rect 433036 291218 433038 291454
rect 432798 291134 433038 291218
rect 432798 290898 432800 291134
rect 433036 290898 433038 291134
rect 432798 290866 433038 290898
rect 433644 291454 433884 291486
rect 433644 291218 433646 291454
rect 433882 291218 433884 291454
rect 433644 291134 433884 291218
rect 433644 290898 433646 291134
rect 433882 290898 433884 291134
rect 433644 290866 433884 290898
rect 442644 291454 442884 291486
rect 442644 291218 442646 291454
rect 442882 291218 442884 291454
rect 442644 291134 442884 291218
rect 442644 290898 442646 291134
rect 442882 290898 442884 291134
rect 442644 290866 442884 290898
rect 451644 291454 451884 291486
rect 451644 291218 451646 291454
rect 451882 291218 451884 291454
rect 451644 291134 451884 291218
rect 451644 290898 451646 291134
rect 451882 290898 451884 291134
rect 451644 290866 451884 290898
rect 460644 291454 460884 291486
rect 460644 291218 460646 291454
rect 460882 291218 460884 291454
rect 460644 291134 460884 291218
rect 460644 290898 460646 291134
rect 460882 290898 460884 291134
rect 460644 290866 460884 290898
rect 469644 291454 469884 291486
rect 469644 291218 469646 291454
rect 469882 291218 469884 291454
rect 469644 291134 469884 291218
rect 469644 290898 469646 291134
rect 469882 290898 469884 291134
rect 469644 290866 469884 290898
rect 471446 291454 471686 291486
rect 471446 291218 471448 291454
rect 471684 291218 471686 291454
rect 471446 291134 471686 291218
rect 471446 290898 471448 291134
rect 471684 290898 471686 291134
rect 471446 290866 471686 290898
rect 578488 291454 579088 291486
rect 578488 291218 578670 291454
rect 578906 291218 579088 291454
rect 578488 291134 579088 291218
rect 578488 290898 578670 291134
rect 578906 290898 579088 291134
rect 578488 290866 579088 290898
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 4400 273454 5000 273486
rect 4400 273218 4582 273454
rect 4818 273218 5000 273454
rect 4400 273134 5000 273218
rect 4400 272898 4582 273134
rect 4818 272898 5000 273134
rect 4400 272866 5000 272898
rect 108278 273454 108518 273486
rect 108278 273218 108280 273454
rect 108516 273218 108518 273454
rect 108278 273134 108518 273218
rect 108278 272898 108280 273134
rect 108516 272898 108518 273134
rect 108278 272866 108518 272898
rect 109084 273454 109324 273486
rect 109084 273218 109086 273454
rect 109322 273218 109324 273454
rect 109084 273134 109324 273218
rect 109084 272898 109086 273134
rect 109322 272898 109324 273134
rect 109084 272866 109324 272898
rect 118084 273454 118324 273486
rect 118084 273218 118086 273454
rect 118322 273218 118324 273454
rect 118084 273134 118324 273218
rect 118084 272898 118086 273134
rect 118322 272898 118324 273134
rect 118084 272866 118324 272898
rect 127084 273454 127324 273486
rect 127084 273218 127086 273454
rect 127322 273218 127324 273454
rect 127084 273134 127324 273218
rect 127084 272898 127086 273134
rect 127322 272898 127324 273134
rect 127084 272866 127324 272898
rect 136084 273454 136324 273486
rect 136084 273218 136086 273454
rect 136322 273218 136324 273454
rect 136084 273134 136324 273218
rect 136084 272898 136086 273134
rect 136322 272898 136324 273134
rect 136084 272866 136324 272898
rect 145084 273454 145324 273486
rect 145084 273218 145086 273454
rect 145322 273218 145324 273454
rect 145084 273134 145324 273218
rect 145084 272898 145086 273134
rect 145322 272898 145324 273134
rect 145084 272866 145324 272898
rect 147646 273454 147886 273486
rect 147646 273218 147648 273454
rect 147884 273218 147886 273454
rect 147646 273134 147886 273218
rect 147646 272898 147648 273134
rect 147884 272898 147886 273134
rect 147646 272866 147886 272898
rect 148780 273454 149020 273486
rect 148780 273218 148782 273454
rect 149018 273218 149020 273454
rect 148780 273134 149020 273218
rect 148780 272898 148782 273134
rect 149018 272898 149020 273134
rect 148780 272866 149020 272898
rect 149298 273454 149538 273486
rect 149298 273218 149300 273454
rect 149536 273218 149538 273454
rect 149298 273134 149538 273218
rect 149298 272898 149300 273134
rect 149536 272898 149538 273134
rect 149298 272866 149538 272898
rect 150104 273454 150344 273486
rect 150104 273218 150106 273454
rect 150342 273218 150344 273454
rect 150104 273134 150344 273218
rect 150104 272898 150106 273134
rect 150342 272898 150344 273134
rect 150104 272866 150344 272898
rect 159104 273454 159344 273486
rect 159104 273218 159106 273454
rect 159342 273218 159344 273454
rect 159104 273134 159344 273218
rect 159104 272898 159106 273134
rect 159342 272898 159344 273134
rect 159104 272866 159344 272898
rect 168104 273454 168344 273486
rect 168104 273218 168106 273454
rect 168342 273218 168344 273454
rect 168104 273134 168344 273218
rect 168104 272898 168106 273134
rect 168342 272898 168344 273134
rect 168104 272866 168344 272898
rect 177104 273454 177344 273486
rect 177104 273218 177106 273454
rect 177342 273218 177344 273454
rect 177104 273134 177344 273218
rect 177104 272898 177106 273134
rect 177342 272898 177344 273134
rect 177104 272866 177344 272898
rect 186104 273454 186344 273486
rect 186104 273218 186106 273454
rect 186342 273218 186344 273454
rect 186104 273134 186344 273218
rect 186104 272898 186106 273134
rect 186342 272898 186344 273134
rect 186104 272866 186344 272898
rect 188666 273454 188906 273486
rect 188666 273218 188668 273454
rect 188904 273218 188906 273454
rect 188666 273134 188906 273218
rect 188666 272898 188668 273134
rect 188904 272898 188906 273134
rect 188666 272866 188906 272898
rect 189214 273454 189454 273486
rect 189214 273218 189216 273454
rect 189452 273218 189454 273454
rect 189214 273134 189454 273218
rect 189214 272898 189216 273134
rect 189452 272898 189454 273134
rect 189214 272866 189454 272898
rect 190318 273454 190558 273486
rect 190318 273218 190320 273454
rect 190556 273218 190558 273454
rect 190318 273134 190558 273218
rect 190318 272898 190320 273134
rect 190556 272898 190558 273134
rect 190318 272866 190558 272898
rect 191124 273454 191364 273486
rect 191124 273218 191126 273454
rect 191362 273218 191364 273454
rect 191124 273134 191364 273218
rect 191124 272898 191126 273134
rect 191362 272898 191364 273134
rect 191124 272866 191364 272898
rect 200124 273454 200364 273486
rect 200124 273218 200126 273454
rect 200362 273218 200364 273454
rect 200124 273134 200364 273218
rect 200124 272898 200126 273134
rect 200362 272898 200364 273134
rect 200124 272866 200364 272898
rect 209124 273454 209364 273486
rect 209124 273218 209126 273454
rect 209362 273218 209364 273454
rect 209124 273134 209364 273218
rect 209124 272898 209126 273134
rect 209362 272898 209364 273134
rect 209124 272866 209364 272898
rect 218124 273454 218364 273486
rect 218124 273218 218126 273454
rect 218362 273218 218364 273454
rect 218124 273134 218364 273218
rect 218124 272898 218126 273134
rect 218362 272898 218364 273134
rect 218124 272866 218364 272898
rect 227124 273454 227364 273486
rect 227124 273218 227126 273454
rect 227362 273218 227364 273454
rect 227124 273134 227364 273218
rect 227124 272898 227126 273134
rect 227362 272898 227364 273134
rect 227124 272866 227364 272898
rect 229686 273454 229926 273486
rect 229686 273218 229688 273454
rect 229924 273218 229926 273454
rect 229686 273134 229926 273218
rect 229686 272898 229688 273134
rect 229924 272898 229926 273134
rect 229686 272866 229926 272898
rect 230338 273454 230578 273486
rect 230338 273218 230340 273454
rect 230576 273218 230578 273454
rect 230338 273134 230578 273218
rect 230338 272898 230340 273134
rect 230576 272898 230578 273134
rect 230338 272866 230578 272898
rect 231144 273454 231384 273486
rect 231144 273218 231146 273454
rect 231382 273218 231384 273454
rect 231144 273134 231384 273218
rect 231144 272898 231146 273134
rect 231382 272898 231384 273134
rect 231144 272866 231384 272898
rect 240144 273454 240384 273486
rect 240144 273218 240146 273454
rect 240382 273218 240384 273454
rect 240144 273134 240384 273218
rect 240144 272898 240146 273134
rect 240382 272898 240384 273134
rect 240144 272866 240384 272898
rect 249144 273454 249384 273486
rect 249144 273218 249146 273454
rect 249382 273218 249384 273454
rect 249144 273134 249384 273218
rect 249144 272898 249146 273134
rect 249382 272898 249384 273134
rect 249144 272866 249384 272898
rect 258144 273454 258384 273486
rect 258144 273218 258146 273454
rect 258382 273218 258384 273454
rect 258144 273134 258384 273218
rect 258144 272898 258146 273134
rect 258382 272898 258384 273134
rect 258144 272866 258384 272898
rect 267144 273454 267384 273486
rect 267144 273218 267146 273454
rect 267382 273218 267384 273454
rect 267144 273134 267384 273218
rect 267144 272898 267146 273134
rect 267382 272898 267384 273134
rect 267144 272866 267384 272898
rect 269706 273454 269946 273486
rect 269706 273218 269708 273454
rect 269944 273218 269946 273454
rect 269706 273134 269946 273218
rect 269706 272898 269708 273134
rect 269944 272898 269946 273134
rect 269706 272866 269946 272898
rect 270358 273454 270598 273486
rect 270358 273218 270360 273454
rect 270596 273218 270598 273454
rect 270358 273134 270598 273218
rect 270358 272898 270360 273134
rect 270596 272898 270598 273134
rect 270358 272866 270598 272898
rect 271164 273454 271404 273486
rect 271164 273218 271166 273454
rect 271402 273218 271404 273454
rect 271164 273134 271404 273218
rect 271164 272898 271166 273134
rect 271402 272898 271404 273134
rect 271164 272866 271404 272898
rect 280164 273454 280404 273486
rect 280164 273218 280166 273454
rect 280402 273218 280404 273454
rect 280164 273134 280404 273218
rect 280164 272898 280166 273134
rect 280402 272898 280404 273134
rect 280164 272866 280404 272898
rect 289164 273454 289404 273486
rect 289164 273218 289166 273454
rect 289402 273218 289404 273454
rect 289164 273134 289404 273218
rect 289164 272898 289166 273134
rect 289402 272898 289404 273134
rect 289164 272866 289404 272898
rect 298164 273454 298404 273486
rect 298164 273218 298166 273454
rect 298402 273218 298404 273454
rect 298164 273134 298404 273218
rect 298164 272898 298166 273134
rect 298402 272898 298404 273134
rect 298164 272866 298404 272898
rect 307164 273454 307404 273486
rect 307164 273218 307166 273454
rect 307402 273218 307404 273454
rect 307164 273134 307404 273218
rect 307164 272898 307166 273134
rect 307402 272898 307404 273134
rect 307164 272866 307404 272898
rect 309726 273454 309966 273486
rect 309726 273218 309728 273454
rect 309964 273218 309966 273454
rect 309726 273134 309966 273218
rect 309726 272898 309728 273134
rect 309964 272898 309966 273134
rect 309726 272866 309966 272898
rect 310838 273454 311078 273486
rect 310838 273218 310840 273454
rect 311076 273218 311078 273454
rect 310838 273134 311078 273218
rect 310838 272898 310840 273134
rect 311076 272898 311078 273134
rect 310838 272866 311078 272898
rect 311378 273454 311618 273486
rect 311378 273218 311380 273454
rect 311616 273218 311618 273454
rect 311378 273134 311618 273218
rect 311378 272898 311380 273134
rect 311616 272898 311618 273134
rect 311378 272866 311618 272898
rect 312184 273454 312424 273486
rect 312184 273218 312186 273454
rect 312422 273218 312424 273454
rect 312184 273134 312424 273218
rect 312184 272898 312186 273134
rect 312422 272898 312424 273134
rect 312184 272866 312424 272898
rect 321184 273454 321424 273486
rect 321184 273218 321186 273454
rect 321422 273218 321424 273454
rect 321184 273134 321424 273218
rect 321184 272898 321186 273134
rect 321422 272898 321424 273134
rect 321184 272866 321424 272898
rect 330184 273454 330424 273486
rect 330184 273218 330186 273454
rect 330422 273218 330424 273454
rect 330184 273134 330424 273218
rect 330184 272898 330186 273134
rect 330422 272898 330424 273134
rect 330184 272866 330424 272898
rect 339184 273454 339424 273486
rect 339184 273218 339186 273454
rect 339422 273218 339424 273454
rect 339184 273134 339424 273218
rect 339184 272898 339186 273134
rect 339422 272898 339424 273134
rect 339184 272866 339424 272898
rect 348184 273454 348424 273486
rect 348184 273218 348186 273454
rect 348422 273218 348424 273454
rect 348184 273134 348424 273218
rect 348184 272898 348186 273134
rect 348422 272898 348424 273134
rect 348184 272866 348424 272898
rect 350746 273454 350986 273486
rect 350746 273218 350748 273454
rect 350984 273218 350986 273454
rect 350746 273134 350986 273218
rect 350746 272898 350748 273134
rect 350984 272898 350986 273134
rect 350746 272866 350986 272898
rect 351318 273454 351558 273486
rect 351318 273218 351320 273454
rect 351556 273218 351558 273454
rect 351318 273134 351558 273218
rect 351318 272898 351320 273134
rect 351556 272898 351558 273134
rect 351318 272866 351558 272898
rect 352398 273454 352638 273486
rect 352398 273218 352400 273454
rect 352636 273218 352638 273454
rect 352398 273134 352638 273218
rect 352398 272898 352400 273134
rect 352636 272898 352638 273134
rect 352398 272866 352638 272898
rect 353204 273454 353444 273486
rect 353204 273218 353206 273454
rect 353442 273218 353444 273454
rect 353204 273134 353444 273218
rect 353204 272898 353206 273134
rect 353442 272898 353444 273134
rect 353204 272866 353444 272898
rect 362204 273454 362444 273486
rect 362204 273218 362206 273454
rect 362442 273218 362444 273454
rect 362204 273134 362444 273218
rect 362204 272898 362206 273134
rect 362442 272898 362444 273134
rect 362204 272866 362444 272898
rect 371204 273454 371444 273486
rect 371204 273218 371206 273454
rect 371442 273218 371444 273454
rect 371204 273134 371444 273218
rect 371204 272898 371206 273134
rect 371442 272898 371444 273134
rect 371204 272866 371444 272898
rect 380204 273454 380444 273486
rect 380204 273218 380206 273454
rect 380442 273218 380444 273454
rect 380204 273134 380444 273218
rect 380204 272898 380206 273134
rect 380442 272898 380444 273134
rect 380204 272866 380444 272898
rect 389204 273454 389444 273486
rect 389204 273218 389206 273454
rect 389442 273218 389444 273454
rect 389204 273134 389444 273218
rect 389204 272898 389206 273134
rect 389442 272898 389444 273134
rect 389204 272866 389444 272898
rect 391766 273454 392006 273486
rect 391766 273218 391768 273454
rect 392004 273218 392006 273454
rect 391766 273134 392006 273218
rect 391766 272898 391768 273134
rect 392004 272898 392006 273134
rect 391766 272866 392006 272898
rect 392418 273454 392658 273486
rect 392418 273218 392420 273454
rect 392656 273218 392658 273454
rect 392418 273134 392658 273218
rect 392418 272898 392420 273134
rect 392656 272898 392658 273134
rect 392418 272866 392658 272898
rect 393224 273454 393464 273486
rect 393224 273218 393226 273454
rect 393462 273218 393464 273454
rect 393224 273134 393464 273218
rect 393224 272898 393226 273134
rect 393462 272898 393464 273134
rect 393224 272866 393464 272898
rect 402224 273454 402464 273486
rect 402224 273218 402226 273454
rect 402462 273218 402464 273454
rect 402224 273134 402464 273218
rect 402224 272898 402226 273134
rect 402462 272898 402464 273134
rect 402224 272866 402464 272898
rect 411224 273454 411464 273486
rect 411224 273218 411226 273454
rect 411462 273218 411464 273454
rect 411224 273134 411464 273218
rect 411224 272898 411226 273134
rect 411462 272898 411464 273134
rect 411224 272866 411464 272898
rect 420224 273454 420464 273486
rect 420224 273218 420226 273454
rect 420462 273218 420464 273454
rect 420224 273134 420464 273218
rect 420224 272898 420226 273134
rect 420462 272898 420464 273134
rect 420224 272866 420464 272898
rect 429224 273454 429464 273486
rect 429224 273218 429226 273454
rect 429462 273218 429464 273454
rect 429224 273134 429464 273218
rect 429224 272898 429226 273134
rect 429462 272898 429464 273134
rect 429224 272866 429464 272898
rect 431786 273454 432026 273486
rect 431786 273218 431788 273454
rect 432024 273218 432026 273454
rect 431786 273134 432026 273218
rect 431786 272898 431788 273134
rect 432024 272898 432026 273134
rect 431786 272866 432026 272898
rect 432438 273454 432678 273486
rect 432438 273218 432440 273454
rect 432676 273218 432678 273454
rect 432438 273134 432678 273218
rect 432438 272898 432440 273134
rect 432676 272898 432678 273134
rect 432438 272866 432678 272898
rect 433244 273454 433484 273486
rect 433244 273218 433246 273454
rect 433482 273218 433484 273454
rect 433244 273134 433484 273218
rect 433244 272898 433246 273134
rect 433482 272898 433484 273134
rect 433244 272866 433484 272898
rect 442244 273454 442484 273486
rect 442244 273218 442246 273454
rect 442482 273218 442484 273454
rect 442244 273134 442484 273218
rect 442244 272898 442246 273134
rect 442482 272898 442484 273134
rect 442244 272866 442484 272898
rect 451244 273454 451484 273486
rect 451244 273218 451246 273454
rect 451482 273218 451484 273454
rect 451244 273134 451484 273218
rect 451244 272898 451246 273134
rect 451482 272898 451484 273134
rect 451244 272866 451484 272898
rect 460244 273454 460484 273486
rect 460244 273218 460246 273454
rect 460482 273218 460484 273454
rect 460244 273134 460484 273218
rect 460244 272898 460246 273134
rect 460482 272898 460484 273134
rect 460244 272866 460484 272898
rect 469244 273454 469484 273486
rect 469244 273218 469246 273454
rect 469482 273218 469484 273454
rect 469244 273134 469484 273218
rect 469244 272898 469246 273134
rect 469482 272898 469484 273134
rect 469244 272866 469484 272898
rect 471806 273454 472046 273486
rect 471806 273218 471808 273454
rect 472044 273218 472046 273454
rect 471806 273134 472046 273218
rect 471806 272898 471808 273134
rect 472044 272898 472046 273134
rect 471806 272866 472046 272898
rect 579288 273454 579888 273486
rect 579288 273218 579470 273454
rect 579706 273218 579888 273454
rect 579288 273134 579888 273218
rect 579288 272898 579470 273134
rect 579706 272898 579888 273134
rect 579288 272866 579888 272898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect 5200 255454 5800 255486
rect 5200 255218 5382 255454
rect 5618 255218 5800 255454
rect 5200 255134 5800 255218
rect 5200 254898 5382 255134
rect 5618 254898 5800 255134
rect 5200 254866 5800 254898
rect 12590 255454 12830 255486
rect 12590 255218 12592 255454
rect 12828 255218 12830 255454
rect 12590 255134 12830 255218
rect 12590 254898 12592 255134
rect 12828 254898 12830 255134
rect 12590 254866 12830 254898
rect 13436 255454 13676 255486
rect 13436 255218 13438 255454
rect 13674 255218 13676 255454
rect 13436 255134 13676 255218
rect 13436 254898 13438 255134
rect 13674 254898 13676 255134
rect 13436 254866 13676 254898
rect 22436 255454 22676 255486
rect 22436 255218 22438 255454
rect 22674 255218 22676 255454
rect 22436 255134 22676 255218
rect 22436 254898 22438 255134
rect 22674 254898 22676 255134
rect 22436 254866 22676 254898
rect 27226 255454 27466 255486
rect 27226 255218 27228 255454
rect 27464 255218 27466 255454
rect 27226 255134 27466 255218
rect 27226 254898 27228 255134
rect 27464 254898 27466 255134
rect 27226 254866 27466 254898
rect 28598 255454 28838 255486
rect 28598 255218 28600 255454
rect 28836 255218 28838 255454
rect 28598 255134 28838 255218
rect 28598 254898 28600 255134
rect 28836 254898 28838 255134
rect 28598 254866 28838 254898
rect 29444 255454 29684 255486
rect 29444 255218 29446 255454
rect 29682 255218 29684 255454
rect 29444 255134 29684 255218
rect 29444 254898 29446 255134
rect 29682 254898 29684 255134
rect 29444 254866 29684 254898
rect 38444 255454 38684 255486
rect 38444 255218 38446 255454
rect 38682 255218 38684 255454
rect 38444 255134 38684 255218
rect 38444 254898 38446 255134
rect 38682 254898 38684 255134
rect 38444 254866 38684 254898
rect 47444 255454 47684 255486
rect 47444 255218 47446 255454
rect 47682 255218 47684 255454
rect 47444 255134 47684 255218
rect 47444 254898 47446 255134
rect 47682 254898 47684 255134
rect 47444 254866 47684 254898
rect 56444 255454 56684 255486
rect 56444 255218 56446 255454
rect 56682 255218 56684 255454
rect 56444 255134 56684 255218
rect 56444 254898 56446 255134
rect 56682 254898 56684 255134
rect 56444 254866 56684 254898
rect 65444 255454 65684 255486
rect 65444 255218 65446 255454
rect 65682 255218 65684 255454
rect 65444 255134 65684 255218
rect 65444 254898 65446 255134
rect 65682 254898 65684 255134
rect 65444 254866 65684 254898
rect 67246 255454 67486 255486
rect 67246 255218 67248 255454
rect 67484 255218 67486 255454
rect 67246 255134 67486 255218
rect 67246 254898 67248 255134
rect 67484 254898 67486 255134
rect 67246 254866 67486 254898
rect 68618 255454 68858 255486
rect 68618 255218 68620 255454
rect 68856 255218 68858 255454
rect 68618 255134 68858 255218
rect 68618 254898 68620 255134
rect 68856 254898 68858 255134
rect 68618 254866 68858 254898
rect 69464 255454 69704 255486
rect 69464 255218 69466 255454
rect 69702 255218 69704 255454
rect 69464 255134 69704 255218
rect 69464 254898 69466 255134
rect 69702 254898 69704 255134
rect 69464 254866 69704 254898
rect 78464 255454 78704 255486
rect 78464 255218 78466 255454
rect 78702 255218 78704 255454
rect 78464 255134 78704 255218
rect 78464 254898 78466 255134
rect 78702 254898 78704 255134
rect 78464 254866 78704 254898
rect 87464 255454 87704 255486
rect 87464 255218 87466 255454
rect 87702 255218 87704 255454
rect 87464 255134 87704 255218
rect 87464 254898 87466 255134
rect 87702 254898 87704 255134
rect 87464 254866 87704 254898
rect 96464 255454 96704 255486
rect 96464 255218 96466 255454
rect 96702 255218 96704 255454
rect 96464 255134 96704 255218
rect 96464 254898 96466 255134
rect 96702 254898 96704 255134
rect 96464 254866 96704 254898
rect 105464 255454 105704 255486
rect 105464 255218 105466 255454
rect 105702 255218 105704 255454
rect 105464 255134 105704 255218
rect 105464 254898 105466 255134
rect 105702 254898 105704 255134
rect 105464 254866 105704 254898
rect 107266 255454 107506 255486
rect 107266 255218 107268 255454
rect 107504 255218 107506 255454
rect 107266 255134 107506 255218
rect 107266 254898 107268 255134
rect 107504 254898 107506 255134
rect 107266 254866 107506 254898
rect 108638 255454 108878 255486
rect 108638 255218 108640 255454
rect 108876 255218 108878 255454
rect 108638 255134 108878 255218
rect 108638 254898 108640 255134
rect 108876 254898 108878 255134
rect 108638 254866 108878 254898
rect 109484 255454 109724 255486
rect 109484 255218 109486 255454
rect 109722 255218 109724 255454
rect 109484 255134 109724 255218
rect 109484 254898 109486 255134
rect 109722 254898 109724 255134
rect 109484 254866 109724 254898
rect 118484 255454 118724 255486
rect 118484 255218 118486 255454
rect 118722 255218 118724 255454
rect 118484 255134 118724 255218
rect 118484 254898 118486 255134
rect 118722 254898 118724 255134
rect 118484 254866 118724 254898
rect 127484 255454 127724 255486
rect 127484 255218 127486 255454
rect 127722 255218 127724 255454
rect 127484 255134 127724 255218
rect 127484 254898 127486 255134
rect 127722 254898 127724 255134
rect 127484 254866 127724 254898
rect 136484 255454 136724 255486
rect 136484 255218 136486 255454
rect 136722 255218 136724 255454
rect 136484 255134 136724 255218
rect 136484 254898 136486 255134
rect 136722 254898 136724 255134
rect 136484 254866 136724 254898
rect 145484 255454 145724 255486
rect 145484 255218 145486 255454
rect 145722 255218 145724 255454
rect 145484 255134 145724 255218
rect 145484 254898 145486 255134
rect 145722 254898 145724 255134
rect 145484 254866 145724 254898
rect 147286 255454 147526 255486
rect 147286 255218 147288 255454
rect 147524 255218 147526 255454
rect 147286 255134 147526 255218
rect 147286 254898 147288 255134
rect 147524 254898 147526 255134
rect 147286 254866 147526 254898
rect 149658 255454 149898 255486
rect 149658 255218 149660 255454
rect 149896 255218 149898 255454
rect 149658 255134 149898 255218
rect 149658 254898 149660 255134
rect 149896 254898 149898 255134
rect 149658 254866 149898 254898
rect 150504 255454 150744 255486
rect 150504 255218 150506 255454
rect 150742 255218 150744 255454
rect 150504 255134 150744 255218
rect 150504 254898 150506 255134
rect 150742 254898 150744 255134
rect 150504 254866 150744 254898
rect 159504 255454 159744 255486
rect 159504 255218 159506 255454
rect 159742 255218 159744 255454
rect 159504 255134 159744 255218
rect 159504 254898 159506 255134
rect 159742 254898 159744 255134
rect 159504 254866 159744 254898
rect 168504 255454 168744 255486
rect 168504 255218 168506 255454
rect 168742 255218 168744 255454
rect 168504 255134 168744 255218
rect 168504 254898 168506 255134
rect 168742 254898 168744 255134
rect 168504 254866 168744 254898
rect 177504 255454 177744 255486
rect 177504 255218 177506 255454
rect 177742 255218 177744 255454
rect 177504 255134 177744 255218
rect 177504 254898 177506 255134
rect 177742 254898 177744 255134
rect 177504 254866 177744 254898
rect 186504 255454 186744 255486
rect 186504 255218 186506 255454
rect 186742 255218 186744 255454
rect 186504 255134 186744 255218
rect 186504 254898 186506 255134
rect 186742 254898 186744 255134
rect 186504 254866 186744 254898
rect 188306 255454 188546 255486
rect 188306 255218 188308 255454
rect 188544 255218 188546 255454
rect 188306 255134 188546 255218
rect 188306 254898 188308 255134
rect 188544 254898 188546 255134
rect 188306 254866 188546 254898
rect 190678 255454 190918 255486
rect 190678 255218 190680 255454
rect 190916 255218 190918 255454
rect 190678 255134 190918 255218
rect 190678 254898 190680 255134
rect 190916 254898 190918 255134
rect 190678 254866 190918 254898
rect 191524 255454 191764 255486
rect 191524 255218 191526 255454
rect 191762 255218 191764 255454
rect 191524 255134 191764 255218
rect 191524 254898 191526 255134
rect 191762 254898 191764 255134
rect 191524 254866 191764 254898
rect 200524 255454 200764 255486
rect 200524 255218 200526 255454
rect 200762 255218 200764 255454
rect 200524 255134 200764 255218
rect 200524 254898 200526 255134
rect 200762 254898 200764 255134
rect 200524 254866 200764 254898
rect 209524 255454 209764 255486
rect 209524 255218 209526 255454
rect 209762 255218 209764 255454
rect 209524 255134 209764 255218
rect 209524 254898 209526 255134
rect 209762 254898 209764 255134
rect 209524 254866 209764 254898
rect 218524 255454 218764 255486
rect 218524 255218 218526 255454
rect 218762 255218 218764 255454
rect 218524 255134 218764 255218
rect 218524 254898 218526 255134
rect 218762 254898 218764 255134
rect 218524 254866 218764 254898
rect 227524 255454 227764 255486
rect 227524 255218 227526 255454
rect 227762 255218 227764 255454
rect 227524 255134 227764 255218
rect 227524 254898 227526 255134
rect 227762 254898 227764 255134
rect 227524 254866 227764 254898
rect 229326 255454 229566 255486
rect 229326 255218 229328 255454
rect 229564 255218 229566 255454
rect 229326 255134 229566 255218
rect 229326 254898 229328 255134
rect 229564 254898 229566 255134
rect 229326 254866 229566 254898
rect 230698 255454 230938 255486
rect 230698 255218 230700 255454
rect 230936 255218 230938 255454
rect 230698 255134 230938 255218
rect 230698 254898 230700 255134
rect 230936 254898 230938 255134
rect 230698 254866 230938 254898
rect 231544 255454 231784 255486
rect 231544 255218 231546 255454
rect 231782 255218 231784 255454
rect 231544 255134 231784 255218
rect 231544 254898 231546 255134
rect 231782 254898 231784 255134
rect 231544 254866 231784 254898
rect 240544 255454 240784 255486
rect 240544 255218 240546 255454
rect 240782 255218 240784 255454
rect 240544 255134 240784 255218
rect 240544 254898 240546 255134
rect 240782 254898 240784 255134
rect 240544 254866 240784 254898
rect 249544 255454 249784 255486
rect 249544 255218 249546 255454
rect 249782 255218 249784 255454
rect 249544 255134 249784 255218
rect 249544 254898 249546 255134
rect 249782 254898 249784 255134
rect 249544 254866 249784 254898
rect 258544 255454 258784 255486
rect 258544 255218 258546 255454
rect 258782 255218 258784 255454
rect 258544 255134 258784 255218
rect 258544 254898 258546 255134
rect 258782 254898 258784 255134
rect 258544 254866 258784 254898
rect 267544 255454 267784 255486
rect 267544 255218 267546 255454
rect 267782 255218 267784 255454
rect 267544 255134 267784 255218
rect 267544 254898 267546 255134
rect 267782 254898 267784 255134
rect 267544 254866 267784 254898
rect 269346 255454 269586 255486
rect 269346 255218 269348 255454
rect 269584 255218 269586 255454
rect 269346 255134 269586 255218
rect 269346 254898 269348 255134
rect 269584 254898 269586 255134
rect 269346 254866 269586 254898
rect 270718 255454 270958 255486
rect 270718 255218 270720 255454
rect 270956 255218 270958 255454
rect 270718 255134 270958 255218
rect 270718 254898 270720 255134
rect 270956 254898 270958 255134
rect 270718 254866 270958 254898
rect 271564 255454 271804 255486
rect 271564 255218 271566 255454
rect 271802 255218 271804 255454
rect 271564 255134 271804 255218
rect 271564 254898 271566 255134
rect 271802 254898 271804 255134
rect 271564 254866 271804 254898
rect 280564 255454 280804 255486
rect 280564 255218 280566 255454
rect 280802 255218 280804 255454
rect 280564 255134 280804 255218
rect 280564 254898 280566 255134
rect 280802 254898 280804 255134
rect 280564 254866 280804 254898
rect 289564 255454 289804 255486
rect 289564 255218 289566 255454
rect 289802 255218 289804 255454
rect 289564 255134 289804 255218
rect 289564 254898 289566 255134
rect 289802 254898 289804 255134
rect 289564 254866 289804 254898
rect 298564 255454 298804 255486
rect 298564 255218 298566 255454
rect 298802 255218 298804 255454
rect 298564 255134 298804 255218
rect 298564 254898 298566 255134
rect 298802 254898 298804 255134
rect 298564 254866 298804 254898
rect 307564 255454 307804 255486
rect 307564 255218 307566 255454
rect 307802 255218 307804 255454
rect 307564 255134 307804 255218
rect 307564 254898 307566 255134
rect 307802 254898 307804 255134
rect 307564 254866 307804 254898
rect 309366 255454 309606 255486
rect 309366 255218 309368 255454
rect 309604 255218 309606 255454
rect 309366 255134 309606 255218
rect 309366 254898 309368 255134
rect 309604 254898 309606 255134
rect 309366 254866 309606 254898
rect 311738 255454 311978 255486
rect 311738 255218 311740 255454
rect 311976 255218 311978 255454
rect 311738 255134 311978 255218
rect 311738 254898 311740 255134
rect 311976 254898 311978 255134
rect 311738 254866 311978 254898
rect 312584 255454 312824 255486
rect 312584 255218 312586 255454
rect 312822 255218 312824 255454
rect 312584 255134 312824 255218
rect 312584 254898 312586 255134
rect 312822 254898 312824 255134
rect 312584 254866 312824 254898
rect 321584 255454 321824 255486
rect 321584 255218 321586 255454
rect 321822 255218 321824 255454
rect 321584 255134 321824 255218
rect 321584 254898 321586 255134
rect 321822 254898 321824 255134
rect 321584 254866 321824 254898
rect 330584 255454 330824 255486
rect 330584 255218 330586 255454
rect 330822 255218 330824 255454
rect 330584 255134 330824 255218
rect 330584 254898 330586 255134
rect 330822 254898 330824 255134
rect 330584 254866 330824 254898
rect 339584 255454 339824 255486
rect 339584 255218 339586 255454
rect 339822 255218 339824 255454
rect 339584 255134 339824 255218
rect 339584 254898 339586 255134
rect 339822 254898 339824 255134
rect 339584 254866 339824 254898
rect 348584 255454 348824 255486
rect 348584 255218 348586 255454
rect 348822 255218 348824 255454
rect 348584 255134 348824 255218
rect 348584 254898 348586 255134
rect 348822 254898 348824 255134
rect 348584 254866 348824 254898
rect 350386 255454 350626 255486
rect 350386 255218 350388 255454
rect 350624 255218 350626 255454
rect 350386 255134 350626 255218
rect 350386 254898 350388 255134
rect 350624 254898 350626 255134
rect 350386 254866 350626 254898
rect 352758 255454 352998 255486
rect 352758 255218 352760 255454
rect 352996 255218 352998 255454
rect 352758 255134 352998 255218
rect 352758 254898 352760 255134
rect 352996 254898 352998 255134
rect 352758 254866 352998 254898
rect 353604 255454 353844 255486
rect 353604 255218 353606 255454
rect 353842 255218 353844 255454
rect 353604 255134 353844 255218
rect 353604 254898 353606 255134
rect 353842 254898 353844 255134
rect 353604 254866 353844 254898
rect 362604 255454 362844 255486
rect 362604 255218 362606 255454
rect 362842 255218 362844 255454
rect 362604 255134 362844 255218
rect 362604 254898 362606 255134
rect 362842 254898 362844 255134
rect 362604 254866 362844 254898
rect 371604 255454 371844 255486
rect 371604 255218 371606 255454
rect 371842 255218 371844 255454
rect 371604 255134 371844 255218
rect 371604 254898 371606 255134
rect 371842 254898 371844 255134
rect 371604 254866 371844 254898
rect 380604 255454 380844 255486
rect 380604 255218 380606 255454
rect 380842 255218 380844 255454
rect 380604 255134 380844 255218
rect 380604 254898 380606 255134
rect 380842 254898 380844 255134
rect 380604 254866 380844 254898
rect 389604 255454 389844 255486
rect 389604 255218 389606 255454
rect 389842 255218 389844 255454
rect 389604 255134 389844 255218
rect 389604 254898 389606 255134
rect 389842 254898 389844 255134
rect 389604 254866 389844 254898
rect 391406 255454 391646 255486
rect 391406 255218 391408 255454
rect 391644 255218 391646 255454
rect 391406 255134 391646 255218
rect 391406 254898 391408 255134
rect 391644 254898 391646 255134
rect 391406 254866 391646 254898
rect 392778 255454 393018 255486
rect 392778 255218 392780 255454
rect 393016 255218 393018 255454
rect 392778 255134 393018 255218
rect 392778 254898 392780 255134
rect 393016 254898 393018 255134
rect 392778 254866 393018 254898
rect 393624 255454 393864 255486
rect 393624 255218 393626 255454
rect 393862 255218 393864 255454
rect 393624 255134 393864 255218
rect 393624 254898 393626 255134
rect 393862 254898 393864 255134
rect 393624 254866 393864 254898
rect 402624 255454 402864 255486
rect 402624 255218 402626 255454
rect 402862 255218 402864 255454
rect 402624 255134 402864 255218
rect 402624 254898 402626 255134
rect 402862 254898 402864 255134
rect 402624 254866 402864 254898
rect 411624 255454 411864 255486
rect 411624 255218 411626 255454
rect 411862 255218 411864 255454
rect 411624 255134 411864 255218
rect 411624 254898 411626 255134
rect 411862 254898 411864 255134
rect 411624 254866 411864 254898
rect 420624 255454 420864 255486
rect 420624 255218 420626 255454
rect 420862 255218 420864 255454
rect 420624 255134 420864 255218
rect 420624 254898 420626 255134
rect 420862 254898 420864 255134
rect 420624 254866 420864 254898
rect 429624 255454 429864 255486
rect 429624 255218 429626 255454
rect 429862 255218 429864 255454
rect 429624 255134 429864 255218
rect 429624 254898 429626 255134
rect 429862 254898 429864 255134
rect 429624 254866 429864 254898
rect 431426 255454 431666 255486
rect 431426 255218 431428 255454
rect 431664 255218 431666 255454
rect 431426 255134 431666 255218
rect 431426 254898 431428 255134
rect 431664 254898 431666 255134
rect 431426 254866 431666 254898
rect 432798 255454 433038 255486
rect 432798 255218 432800 255454
rect 433036 255218 433038 255454
rect 432798 255134 433038 255218
rect 432798 254898 432800 255134
rect 433036 254898 433038 255134
rect 432798 254866 433038 254898
rect 433644 255454 433884 255486
rect 433644 255218 433646 255454
rect 433882 255218 433884 255454
rect 433644 255134 433884 255218
rect 433644 254898 433646 255134
rect 433882 254898 433884 255134
rect 433644 254866 433884 254898
rect 442644 255454 442884 255486
rect 442644 255218 442646 255454
rect 442882 255218 442884 255454
rect 442644 255134 442884 255218
rect 442644 254898 442646 255134
rect 442882 254898 442884 255134
rect 442644 254866 442884 254898
rect 451644 255454 451884 255486
rect 451644 255218 451646 255454
rect 451882 255218 451884 255454
rect 451644 255134 451884 255218
rect 451644 254898 451646 255134
rect 451882 254898 451884 255134
rect 451644 254866 451884 254898
rect 460644 255454 460884 255486
rect 460644 255218 460646 255454
rect 460882 255218 460884 255454
rect 460644 255134 460884 255218
rect 460644 254898 460646 255134
rect 460882 254898 460884 255134
rect 460644 254866 460884 254898
rect 469644 255454 469884 255486
rect 469644 255218 469646 255454
rect 469882 255218 469884 255454
rect 469644 255134 469884 255218
rect 469644 254898 469646 255134
rect 469882 254898 469884 255134
rect 469644 254866 469884 254898
rect 471446 255454 471686 255486
rect 471446 255218 471448 255454
rect 471684 255218 471686 255454
rect 471446 255134 471686 255218
rect 471446 254898 471448 255134
rect 471684 254898 471686 255134
rect 471446 254866 471686 254898
rect 472818 255454 473058 255486
rect 472818 255218 472820 255454
rect 473056 255218 473058 255454
rect 472818 255134 473058 255218
rect 472818 254898 472820 255134
rect 473056 254898 473058 255134
rect 472818 254866 473058 254898
rect 473664 255454 473904 255486
rect 473664 255218 473666 255454
rect 473902 255218 473904 255454
rect 473664 255134 473904 255218
rect 473664 254898 473666 255134
rect 473902 254898 473904 255134
rect 473664 254866 473904 254898
rect 482664 255454 482904 255486
rect 482664 255218 482666 255454
rect 482902 255218 482904 255454
rect 482664 255134 482904 255218
rect 482664 254898 482666 255134
rect 482902 254898 482904 255134
rect 482664 254866 482904 254898
rect 491664 255454 491904 255486
rect 491664 255218 491666 255454
rect 491902 255218 491904 255454
rect 491664 255134 491904 255218
rect 491664 254898 491666 255134
rect 491902 254898 491904 255134
rect 491664 254866 491904 254898
rect 500664 255454 500904 255486
rect 500664 255218 500666 255454
rect 500902 255218 500904 255454
rect 500664 255134 500904 255218
rect 500664 254898 500666 255134
rect 500902 254898 500904 255134
rect 500664 254866 500904 254898
rect 509664 255454 509904 255486
rect 509664 255218 509666 255454
rect 509902 255218 509904 255454
rect 509664 255134 509904 255218
rect 509664 254898 509666 255134
rect 509902 254898 509904 255134
rect 509664 254866 509904 254898
rect 511466 255454 511706 255486
rect 511466 255218 511468 255454
rect 511704 255218 511706 255454
rect 511466 255134 511706 255218
rect 511466 254898 511468 255134
rect 511704 254898 511706 255134
rect 511466 254866 511706 254898
rect 512838 255454 513078 255486
rect 512838 255218 512840 255454
rect 513076 255218 513078 255454
rect 512838 255134 513078 255218
rect 512838 254898 512840 255134
rect 513076 254898 513078 255134
rect 512838 254866 513078 254898
rect 513684 255454 513924 255486
rect 513684 255218 513686 255454
rect 513922 255218 513924 255454
rect 513684 255134 513924 255218
rect 513684 254898 513686 255134
rect 513922 254898 513924 255134
rect 513684 254866 513924 254898
rect 522684 255454 522924 255486
rect 522684 255218 522686 255454
rect 522922 255218 522924 255454
rect 522684 255134 522924 255218
rect 522684 254898 522686 255134
rect 522922 254898 522924 255134
rect 522684 254866 522924 254898
rect 531684 255454 531924 255486
rect 531684 255218 531686 255454
rect 531922 255218 531924 255454
rect 531684 255134 531924 255218
rect 531684 254898 531686 255134
rect 531922 254898 531924 255134
rect 531684 254866 531924 254898
rect 540684 255454 540924 255486
rect 540684 255218 540686 255454
rect 540922 255218 540924 255454
rect 540684 255134 540924 255218
rect 540684 254898 540686 255134
rect 540922 254898 540924 255134
rect 540684 254866 540924 254898
rect 549684 255454 549924 255486
rect 549684 255218 549686 255454
rect 549922 255218 549924 255454
rect 549684 255134 549924 255218
rect 549684 254898 549686 255134
rect 549922 254898 549924 255134
rect 549684 254866 549924 254898
rect 551486 255454 551726 255486
rect 551486 255218 551488 255454
rect 551724 255218 551726 255454
rect 551486 255134 551726 255218
rect 551486 254898 551488 255134
rect 551724 254898 551726 255134
rect 551486 254866 551726 254898
rect 552858 255454 553098 255486
rect 552858 255218 552860 255454
rect 553096 255218 553098 255454
rect 552858 255134 553098 255218
rect 552858 254898 552860 255134
rect 553096 254898 553098 255134
rect 552858 254866 553098 254898
rect 553704 255454 553944 255486
rect 553704 255218 553706 255454
rect 553942 255218 553944 255454
rect 553704 255134 553944 255218
rect 553704 254898 553706 255134
rect 553942 254898 553944 255134
rect 553704 254866 553944 254898
rect 562704 255454 562944 255486
rect 562704 255218 562706 255454
rect 562942 255218 562944 255454
rect 562704 255134 562944 255218
rect 562704 254898 562706 255134
rect 562942 254898 562944 255134
rect 562704 254866 562944 254898
rect 571704 255454 571944 255486
rect 571704 255218 571706 255454
rect 571942 255218 571944 255454
rect 571704 255134 571944 255218
rect 571704 254898 571706 255134
rect 571942 254898 571944 255134
rect 571704 254866 571944 254898
rect 573474 255454 573714 255486
rect 573474 255218 573476 255454
rect 573712 255218 573714 255454
rect 573474 255134 573714 255218
rect 573474 254898 573476 255134
rect 573712 254898 573714 255134
rect 573474 254866 573714 254898
rect 578488 255454 579088 255486
rect 578488 255218 578670 255454
rect 578906 255218 579088 255454
rect 578488 255134 579088 255218
rect 578488 254898 578670 255134
rect 578906 254898 579088 255134
rect 578488 254866 579088 254898
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 4400 237454 5000 237486
rect 4400 237218 4582 237454
rect 4818 237218 5000 237454
rect 4400 237134 5000 237218
rect 4400 236898 4582 237134
rect 4818 236898 5000 237134
rect 4400 236866 5000 236898
rect 12230 237454 12470 237486
rect 12230 237218 12232 237454
rect 12468 237218 12470 237454
rect 12230 237134 12470 237218
rect 12230 236898 12232 237134
rect 12468 236898 12470 237134
rect 12230 236866 12470 236898
rect 13036 237454 13276 237486
rect 13036 237218 13038 237454
rect 13274 237218 13276 237454
rect 13036 237134 13276 237218
rect 13036 236898 13038 237134
rect 13274 236898 13276 237134
rect 13036 236866 13276 236898
rect 22036 237454 22276 237486
rect 22036 237218 22038 237454
rect 22274 237218 22276 237454
rect 22036 237134 22276 237218
rect 22036 236898 22038 237134
rect 22274 236898 22276 237134
rect 22036 236866 22276 236898
rect 27586 237454 27826 237486
rect 27586 237218 27588 237454
rect 27824 237218 27826 237454
rect 27586 237134 27826 237218
rect 27586 236898 27588 237134
rect 27824 236898 27826 237134
rect 27586 236866 27826 236898
rect 28238 237454 28478 237486
rect 28238 237218 28240 237454
rect 28476 237218 28478 237454
rect 28238 237134 28478 237218
rect 28238 236898 28240 237134
rect 28476 236898 28478 237134
rect 28238 236866 28478 236898
rect 29044 237454 29284 237486
rect 29044 237218 29046 237454
rect 29282 237218 29284 237454
rect 29044 237134 29284 237218
rect 29044 236898 29046 237134
rect 29282 236898 29284 237134
rect 29044 236866 29284 236898
rect 38044 237454 38284 237486
rect 38044 237218 38046 237454
rect 38282 237218 38284 237454
rect 38044 237134 38284 237218
rect 38044 236898 38046 237134
rect 38282 236898 38284 237134
rect 38044 236866 38284 236898
rect 47044 237454 47284 237486
rect 47044 237218 47046 237454
rect 47282 237218 47284 237454
rect 47044 237134 47284 237218
rect 47044 236898 47046 237134
rect 47282 236898 47284 237134
rect 47044 236866 47284 236898
rect 56044 237454 56284 237486
rect 56044 237218 56046 237454
rect 56282 237218 56284 237454
rect 56044 237134 56284 237218
rect 56044 236898 56046 237134
rect 56282 236898 56284 237134
rect 56044 236866 56284 236898
rect 65044 237454 65284 237486
rect 65044 237218 65046 237454
rect 65282 237218 65284 237454
rect 65044 237134 65284 237218
rect 65044 236898 65046 237134
rect 65282 236898 65284 237134
rect 65044 236866 65284 236898
rect 67606 237454 67846 237486
rect 67606 237218 67608 237454
rect 67844 237218 67846 237454
rect 67606 237134 67846 237218
rect 67606 236898 67608 237134
rect 67844 236898 67846 237134
rect 67606 236866 67846 236898
rect 68258 237454 68498 237486
rect 68258 237218 68260 237454
rect 68496 237218 68498 237454
rect 68258 237134 68498 237218
rect 68258 236898 68260 237134
rect 68496 236898 68498 237134
rect 68258 236866 68498 236898
rect 69064 237454 69304 237486
rect 69064 237218 69066 237454
rect 69302 237218 69304 237454
rect 69064 237134 69304 237218
rect 69064 236898 69066 237134
rect 69302 236898 69304 237134
rect 69064 236866 69304 236898
rect 78064 237454 78304 237486
rect 78064 237218 78066 237454
rect 78302 237218 78304 237454
rect 78064 237134 78304 237218
rect 78064 236898 78066 237134
rect 78302 236898 78304 237134
rect 78064 236866 78304 236898
rect 87064 237454 87304 237486
rect 87064 237218 87066 237454
rect 87302 237218 87304 237454
rect 87064 237134 87304 237218
rect 87064 236898 87066 237134
rect 87302 236898 87304 237134
rect 87064 236866 87304 236898
rect 96064 237454 96304 237486
rect 96064 237218 96066 237454
rect 96302 237218 96304 237454
rect 96064 237134 96304 237218
rect 96064 236898 96066 237134
rect 96302 236898 96304 237134
rect 96064 236866 96304 236898
rect 105064 237454 105304 237486
rect 105064 237218 105066 237454
rect 105302 237218 105304 237454
rect 105064 237134 105304 237218
rect 105064 236898 105066 237134
rect 105302 236898 105304 237134
rect 105064 236866 105304 236898
rect 107626 237454 107866 237486
rect 107626 237218 107628 237454
rect 107864 237218 107866 237454
rect 107626 237134 107866 237218
rect 107626 236898 107628 237134
rect 107864 236898 107866 237134
rect 107626 236866 107866 236898
rect 108278 237454 108518 237486
rect 108278 237218 108280 237454
rect 108516 237218 108518 237454
rect 108278 237134 108518 237218
rect 108278 236898 108280 237134
rect 108516 236898 108518 237134
rect 108278 236866 108518 236898
rect 109084 237454 109324 237486
rect 109084 237218 109086 237454
rect 109322 237218 109324 237454
rect 109084 237134 109324 237218
rect 109084 236898 109086 237134
rect 109322 236898 109324 237134
rect 109084 236866 109324 236898
rect 118084 237454 118324 237486
rect 118084 237218 118086 237454
rect 118322 237218 118324 237454
rect 118084 237134 118324 237218
rect 118084 236898 118086 237134
rect 118322 236898 118324 237134
rect 118084 236866 118324 236898
rect 127084 237454 127324 237486
rect 127084 237218 127086 237454
rect 127322 237218 127324 237454
rect 127084 237134 127324 237218
rect 127084 236898 127086 237134
rect 127322 236898 127324 237134
rect 127084 236866 127324 236898
rect 136084 237454 136324 237486
rect 136084 237218 136086 237454
rect 136322 237218 136324 237454
rect 136084 237134 136324 237218
rect 136084 236898 136086 237134
rect 136322 236898 136324 237134
rect 136084 236866 136324 236898
rect 145084 237454 145324 237486
rect 145084 237218 145086 237454
rect 145322 237218 145324 237454
rect 145084 237134 145324 237218
rect 145084 236898 145086 237134
rect 145322 236898 145324 237134
rect 145084 236866 145324 236898
rect 147646 237454 147886 237486
rect 147646 237218 147648 237454
rect 147884 237218 147886 237454
rect 147646 237134 147886 237218
rect 147646 236898 147648 237134
rect 147884 236898 147886 237134
rect 147646 236866 147886 236898
rect 148780 237454 149020 237486
rect 148780 237218 148782 237454
rect 149018 237218 149020 237454
rect 148780 237134 149020 237218
rect 148780 236898 148782 237134
rect 149018 236898 149020 237134
rect 148780 236866 149020 236898
rect 149298 237454 149538 237486
rect 149298 237218 149300 237454
rect 149536 237218 149538 237454
rect 149298 237134 149538 237218
rect 149298 236898 149300 237134
rect 149536 236898 149538 237134
rect 149298 236866 149538 236898
rect 150104 237454 150344 237486
rect 150104 237218 150106 237454
rect 150342 237218 150344 237454
rect 150104 237134 150344 237218
rect 150104 236898 150106 237134
rect 150342 236898 150344 237134
rect 150104 236866 150344 236898
rect 159104 237454 159344 237486
rect 159104 237218 159106 237454
rect 159342 237218 159344 237454
rect 159104 237134 159344 237218
rect 159104 236898 159106 237134
rect 159342 236898 159344 237134
rect 159104 236866 159344 236898
rect 168104 237454 168344 237486
rect 168104 237218 168106 237454
rect 168342 237218 168344 237454
rect 168104 237134 168344 237218
rect 168104 236898 168106 237134
rect 168342 236898 168344 237134
rect 168104 236866 168344 236898
rect 177104 237454 177344 237486
rect 177104 237218 177106 237454
rect 177342 237218 177344 237454
rect 177104 237134 177344 237218
rect 177104 236898 177106 237134
rect 177342 236898 177344 237134
rect 177104 236866 177344 236898
rect 186104 237454 186344 237486
rect 186104 237218 186106 237454
rect 186342 237218 186344 237454
rect 186104 237134 186344 237218
rect 186104 236898 186106 237134
rect 186342 236898 186344 237134
rect 186104 236866 186344 236898
rect 188666 237454 188906 237486
rect 188666 237218 188668 237454
rect 188904 237218 188906 237454
rect 188666 237134 188906 237218
rect 188666 236898 188668 237134
rect 188904 236898 188906 237134
rect 188666 236866 188906 236898
rect 189214 237454 189454 237486
rect 189214 237218 189216 237454
rect 189452 237218 189454 237454
rect 189214 237134 189454 237218
rect 189214 236898 189216 237134
rect 189452 236898 189454 237134
rect 189214 236866 189454 236898
rect 190318 237454 190558 237486
rect 190318 237218 190320 237454
rect 190556 237218 190558 237454
rect 190318 237134 190558 237218
rect 190318 236898 190320 237134
rect 190556 236898 190558 237134
rect 190318 236866 190558 236898
rect 191124 237454 191364 237486
rect 191124 237218 191126 237454
rect 191362 237218 191364 237454
rect 191124 237134 191364 237218
rect 191124 236898 191126 237134
rect 191362 236898 191364 237134
rect 191124 236866 191364 236898
rect 200124 237454 200364 237486
rect 200124 237218 200126 237454
rect 200362 237218 200364 237454
rect 200124 237134 200364 237218
rect 200124 236898 200126 237134
rect 200362 236898 200364 237134
rect 200124 236866 200364 236898
rect 209124 237454 209364 237486
rect 209124 237218 209126 237454
rect 209362 237218 209364 237454
rect 209124 237134 209364 237218
rect 209124 236898 209126 237134
rect 209362 236898 209364 237134
rect 209124 236866 209364 236898
rect 218124 237454 218364 237486
rect 218124 237218 218126 237454
rect 218362 237218 218364 237454
rect 218124 237134 218364 237218
rect 218124 236898 218126 237134
rect 218362 236898 218364 237134
rect 218124 236866 218364 236898
rect 227124 237454 227364 237486
rect 227124 237218 227126 237454
rect 227362 237218 227364 237454
rect 227124 237134 227364 237218
rect 227124 236898 227126 237134
rect 227362 236898 227364 237134
rect 227124 236866 227364 236898
rect 229686 237454 229926 237486
rect 229686 237218 229688 237454
rect 229924 237218 229926 237454
rect 229686 237134 229926 237218
rect 229686 236898 229688 237134
rect 229924 236898 229926 237134
rect 229686 236866 229926 236898
rect 230338 237454 230578 237486
rect 230338 237218 230340 237454
rect 230576 237218 230578 237454
rect 230338 237134 230578 237218
rect 230338 236898 230340 237134
rect 230576 236898 230578 237134
rect 230338 236866 230578 236898
rect 231144 237454 231384 237486
rect 231144 237218 231146 237454
rect 231382 237218 231384 237454
rect 231144 237134 231384 237218
rect 231144 236898 231146 237134
rect 231382 236898 231384 237134
rect 231144 236866 231384 236898
rect 240144 237454 240384 237486
rect 240144 237218 240146 237454
rect 240382 237218 240384 237454
rect 240144 237134 240384 237218
rect 240144 236898 240146 237134
rect 240382 236898 240384 237134
rect 240144 236866 240384 236898
rect 249144 237454 249384 237486
rect 249144 237218 249146 237454
rect 249382 237218 249384 237454
rect 249144 237134 249384 237218
rect 249144 236898 249146 237134
rect 249382 236898 249384 237134
rect 249144 236866 249384 236898
rect 258144 237454 258384 237486
rect 258144 237218 258146 237454
rect 258382 237218 258384 237454
rect 258144 237134 258384 237218
rect 258144 236898 258146 237134
rect 258382 236898 258384 237134
rect 258144 236866 258384 236898
rect 267144 237454 267384 237486
rect 267144 237218 267146 237454
rect 267382 237218 267384 237454
rect 267144 237134 267384 237218
rect 267144 236898 267146 237134
rect 267382 236898 267384 237134
rect 267144 236866 267384 236898
rect 269706 237454 269946 237486
rect 269706 237218 269708 237454
rect 269944 237218 269946 237454
rect 269706 237134 269946 237218
rect 269706 236898 269708 237134
rect 269944 236898 269946 237134
rect 269706 236866 269946 236898
rect 270358 237454 270598 237486
rect 270358 237218 270360 237454
rect 270596 237218 270598 237454
rect 270358 237134 270598 237218
rect 270358 236898 270360 237134
rect 270596 236898 270598 237134
rect 270358 236866 270598 236898
rect 271164 237454 271404 237486
rect 271164 237218 271166 237454
rect 271402 237218 271404 237454
rect 271164 237134 271404 237218
rect 271164 236898 271166 237134
rect 271402 236898 271404 237134
rect 271164 236866 271404 236898
rect 280164 237454 280404 237486
rect 280164 237218 280166 237454
rect 280402 237218 280404 237454
rect 280164 237134 280404 237218
rect 280164 236898 280166 237134
rect 280402 236898 280404 237134
rect 280164 236866 280404 236898
rect 289164 237454 289404 237486
rect 289164 237218 289166 237454
rect 289402 237218 289404 237454
rect 289164 237134 289404 237218
rect 289164 236898 289166 237134
rect 289402 236898 289404 237134
rect 289164 236866 289404 236898
rect 298164 237454 298404 237486
rect 298164 237218 298166 237454
rect 298402 237218 298404 237454
rect 298164 237134 298404 237218
rect 298164 236898 298166 237134
rect 298402 236898 298404 237134
rect 298164 236866 298404 236898
rect 307164 237454 307404 237486
rect 307164 237218 307166 237454
rect 307402 237218 307404 237454
rect 307164 237134 307404 237218
rect 307164 236898 307166 237134
rect 307402 236898 307404 237134
rect 307164 236866 307404 236898
rect 309726 237454 309966 237486
rect 309726 237218 309728 237454
rect 309964 237218 309966 237454
rect 309726 237134 309966 237218
rect 309726 236898 309728 237134
rect 309964 236898 309966 237134
rect 309726 236866 309966 236898
rect 310838 237454 311078 237486
rect 310838 237218 310840 237454
rect 311076 237218 311078 237454
rect 310838 237134 311078 237218
rect 310838 236898 310840 237134
rect 311076 236898 311078 237134
rect 310838 236866 311078 236898
rect 311378 237454 311618 237486
rect 311378 237218 311380 237454
rect 311616 237218 311618 237454
rect 311378 237134 311618 237218
rect 311378 236898 311380 237134
rect 311616 236898 311618 237134
rect 311378 236866 311618 236898
rect 312184 237454 312424 237486
rect 312184 237218 312186 237454
rect 312422 237218 312424 237454
rect 312184 237134 312424 237218
rect 312184 236898 312186 237134
rect 312422 236898 312424 237134
rect 312184 236866 312424 236898
rect 321184 237454 321424 237486
rect 321184 237218 321186 237454
rect 321422 237218 321424 237454
rect 321184 237134 321424 237218
rect 321184 236898 321186 237134
rect 321422 236898 321424 237134
rect 321184 236866 321424 236898
rect 330184 237454 330424 237486
rect 330184 237218 330186 237454
rect 330422 237218 330424 237454
rect 330184 237134 330424 237218
rect 330184 236898 330186 237134
rect 330422 236898 330424 237134
rect 330184 236866 330424 236898
rect 339184 237454 339424 237486
rect 339184 237218 339186 237454
rect 339422 237218 339424 237454
rect 339184 237134 339424 237218
rect 339184 236898 339186 237134
rect 339422 236898 339424 237134
rect 339184 236866 339424 236898
rect 348184 237454 348424 237486
rect 348184 237218 348186 237454
rect 348422 237218 348424 237454
rect 348184 237134 348424 237218
rect 348184 236898 348186 237134
rect 348422 236898 348424 237134
rect 348184 236866 348424 236898
rect 350746 237454 350986 237486
rect 350746 237218 350748 237454
rect 350984 237218 350986 237454
rect 350746 237134 350986 237218
rect 350746 236898 350748 237134
rect 350984 236898 350986 237134
rect 350746 236866 350986 236898
rect 351318 237454 351558 237486
rect 351318 237218 351320 237454
rect 351556 237218 351558 237454
rect 351318 237134 351558 237218
rect 351318 236898 351320 237134
rect 351556 236898 351558 237134
rect 351318 236866 351558 236898
rect 352398 237454 352638 237486
rect 352398 237218 352400 237454
rect 352636 237218 352638 237454
rect 352398 237134 352638 237218
rect 352398 236898 352400 237134
rect 352636 236898 352638 237134
rect 352398 236866 352638 236898
rect 353204 237454 353444 237486
rect 353204 237218 353206 237454
rect 353442 237218 353444 237454
rect 353204 237134 353444 237218
rect 353204 236898 353206 237134
rect 353442 236898 353444 237134
rect 353204 236866 353444 236898
rect 362204 237454 362444 237486
rect 362204 237218 362206 237454
rect 362442 237218 362444 237454
rect 362204 237134 362444 237218
rect 362204 236898 362206 237134
rect 362442 236898 362444 237134
rect 362204 236866 362444 236898
rect 371204 237454 371444 237486
rect 371204 237218 371206 237454
rect 371442 237218 371444 237454
rect 371204 237134 371444 237218
rect 371204 236898 371206 237134
rect 371442 236898 371444 237134
rect 371204 236866 371444 236898
rect 380204 237454 380444 237486
rect 380204 237218 380206 237454
rect 380442 237218 380444 237454
rect 380204 237134 380444 237218
rect 380204 236898 380206 237134
rect 380442 236898 380444 237134
rect 380204 236866 380444 236898
rect 389204 237454 389444 237486
rect 389204 237218 389206 237454
rect 389442 237218 389444 237454
rect 389204 237134 389444 237218
rect 389204 236898 389206 237134
rect 389442 236898 389444 237134
rect 389204 236866 389444 236898
rect 391766 237454 392006 237486
rect 391766 237218 391768 237454
rect 392004 237218 392006 237454
rect 391766 237134 392006 237218
rect 391766 236898 391768 237134
rect 392004 236898 392006 237134
rect 391766 236866 392006 236898
rect 392418 237454 392658 237486
rect 392418 237218 392420 237454
rect 392656 237218 392658 237454
rect 392418 237134 392658 237218
rect 392418 236898 392420 237134
rect 392656 236898 392658 237134
rect 392418 236866 392658 236898
rect 393224 237454 393464 237486
rect 393224 237218 393226 237454
rect 393462 237218 393464 237454
rect 393224 237134 393464 237218
rect 393224 236898 393226 237134
rect 393462 236898 393464 237134
rect 393224 236866 393464 236898
rect 402224 237454 402464 237486
rect 402224 237218 402226 237454
rect 402462 237218 402464 237454
rect 402224 237134 402464 237218
rect 402224 236898 402226 237134
rect 402462 236898 402464 237134
rect 402224 236866 402464 236898
rect 411224 237454 411464 237486
rect 411224 237218 411226 237454
rect 411462 237218 411464 237454
rect 411224 237134 411464 237218
rect 411224 236898 411226 237134
rect 411462 236898 411464 237134
rect 411224 236866 411464 236898
rect 420224 237454 420464 237486
rect 420224 237218 420226 237454
rect 420462 237218 420464 237454
rect 420224 237134 420464 237218
rect 420224 236898 420226 237134
rect 420462 236898 420464 237134
rect 420224 236866 420464 236898
rect 429224 237454 429464 237486
rect 429224 237218 429226 237454
rect 429462 237218 429464 237454
rect 429224 237134 429464 237218
rect 429224 236898 429226 237134
rect 429462 236898 429464 237134
rect 429224 236866 429464 236898
rect 431786 237454 432026 237486
rect 431786 237218 431788 237454
rect 432024 237218 432026 237454
rect 431786 237134 432026 237218
rect 431786 236898 431788 237134
rect 432024 236898 432026 237134
rect 431786 236866 432026 236898
rect 432438 237454 432678 237486
rect 432438 237218 432440 237454
rect 432676 237218 432678 237454
rect 432438 237134 432678 237218
rect 432438 236898 432440 237134
rect 432676 236898 432678 237134
rect 432438 236866 432678 236898
rect 433244 237454 433484 237486
rect 433244 237218 433246 237454
rect 433482 237218 433484 237454
rect 433244 237134 433484 237218
rect 433244 236898 433246 237134
rect 433482 236898 433484 237134
rect 433244 236866 433484 236898
rect 442244 237454 442484 237486
rect 442244 237218 442246 237454
rect 442482 237218 442484 237454
rect 442244 237134 442484 237218
rect 442244 236898 442246 237134
rect 442482 236898 442484 237134
rect 442244 236866 442484 236898
rect 451244 237454 451484 237486
rect 451244 237218 451246 237454
rect 451482 237218 451484 237454
rect 451244 237134 451484 237218
rect 451244 236898 451246 237134
rect 451482 236898 451484 237134
rect 451244 236866 451484 236898
rect 460244 237454 460484 237486
rect 460244 237218 460246 237454
rect 460482 237218 460484 237454
rect 460244 237134 460484 237218
rect 460244 236898 460246 237134
rect 460482 236898 460484 237134
rect 460244 236866 460484 236898
rect 469244 237454 469484 237486
rect 469244 237218 469246 237454
rect 469482 237218 469484 237454
rect 469244 237134 469484 237218
rect 469244 236898 469246 237134
rect 469482 236898 469484 237134
rect 469244 236866 469484 236898
rect 471806 237454 472046 237486
rect 471806 237218 471808 237454
rect 472044 237218 472046 237454
rect 471806 237134 472046 237218
rect 471806 236898 471808 237134
rect 472044 236898 472046 237134
rect 471806 236866 472046 236898
rect 472458 237454 472698 237486
rect 472458 237218 472460 237454
rect 472696 237218 472698 237454
rect 472458 237134 472698 237218
rect 472458 236898 472460 237134
rect 472696 236898 472698 237134
rect 472458 236866 472698 236898
rect 473264 237454 473504 237486
rect 473264 237218 473266 237454
rect 473502 237218 473504 237454
rect 473264 237134 473504 237218
rect 473264 236898 473266 237134
rect 473502 236898 473504 237134
rect 473264 236866 473504 236898
rect 482264 237454 482504 237486
rect 482264 237218 482266 237454
rect 482502 237218 482504 237454
rect 482264 237134 482504 237218
rect 482264 236898 482266 237134
rect 482502 236898 482504 237134
rect 482264 236866 482504 236898
rect 491264 237454 491504 237486
rect 491264 237218 491266 237454
rect 491502 237218 491504 237454
rect 491264 237134 491504 237218
rect 491264 236898 491266 237134
rect 491502 236898 491504 237134
rect 491264 236866 491504 236898
rect 500264 237454 500504 237486
rect 500264 237218 500266 237454
rect 500502 237218 500504 237454
rect 500264 237134 500504 237218
rect 500264 236898 500266 237134
rect 500502 236898 500504 237134
rect 500264 236866 500504 236898
rect 509264 237454 509504 237486
rect 509264 237218 509266 237454
rect 509502 237218 509504 237454
rect 509264 237134 509504 237218
rect 509264 236898 509266 237134
rect 509502 236898 509504 237134
rect 509264 236866 509504 236898
rect 511826 237454 512066 237486
rect 511826 237218 511828 237454
rect 512064 237218 512066 237454
rect 511826 237134 512066 237218
rect 511826 236898 511828 237134
rect 512064 236898 512066 237134
rect 511826 236866 512066 236898
rect 512478 237454 512718 237486
rect 512478 237218 512480 237454
rect 512716 237218 512718 237454
rect 512478 237134 512718 237218
rect 512478 236898 512480 237134
rect 512716 236898 512718 237134
rect 512478 236866 512718 236898
rect 513284 237454 513524 237486
rect 513284 237218 513286 237454
rect 513522 237218 513524 237454
rect 513284 237134 513524 237218
rect 513284 236898 513286 237134
rect 513522 236898 513524 237134
rect 513284 236866 513524 236898
rect 522284 237454 522524 237486
rect 522284 237218 522286 237454
rect 522522 237218 522524 237454
rect 522284 237134 522524 237218
rect 522284 236898 522286 237134
rect 522522 236898 522524 237134
rect 522284 236866 522524 236898
rect 531284 237454 531524 237486
rect 531284 237218 531286 237454
rect 531522 237218 531524 237454
rect 531284 237134 531524 237218
rect 531284 236898 531286 237134
rect 531522 236898 531524 237134
rect 531284 236866 531524 236898
rect 540284 237454 540524 237486
rect 540284 237218 540286 237454
rect 540522 237218 540524 237454
rect 540284 237134 540524 237218
rect 540284 236898 540286 237134
rect 540522 236898 540524 237134
rect 540284 236866 540524 236898
rect 549284 237454 549524 237486
rect 549284 237218 549286 237454
rect 549522 237218 549524 237454
rect 549284 237134 549524 237218
rect 549284 236898 549286 237134
rect 549522 236898 549524 237134
rect 549284 236866 549524 236898
rect 551846 237454 552086 237486
rect 551846 237218 551848 237454
rect 552084 237218 552086 237454
rect 551846 237134 552086 237218
rect 551846 236898 551848 237134
rect 552084 236898 552086 237134
rect 551846 236866 552086 236898
rect 552498 237454 552738 237486
rect 552498 237218 552500 237454
rect 552736 237218 552738 237454
rect 552498 237134 552738 237218
rect 552498 236898 552500 237134
rect 552736 236898 552738 237134
rect 552498 236866 552738 236898
rect 553304 237454 553544 237486
rect 553304 237218 553306 237454
rect 553542 237218 553544 237454
rect 553304 237134 553544 237218
rect 553304 236898 553306 237134
rect 553542 236898 553544 237134
rect 553304 236866 553544 236898
rect 562304 237454 562544 237486
rect 562304 237218 562306 237454
rect 562542 237218 562544 237454
rect 562304 237134 562544 237218
rect 562304 236898 562306 237134
rect 562542 236898 562544 237134
rect 562304 236866 562544 236898
rect 571304 237454 571544 237486
rect 571304 237218 571306 237454
rect 571542 237218 571544 237454
rect 571304 237134 571544 237218
rect 571304 236898 571306 237134
rect 571542 236898 571544 237134
rect 571304 236866 571544 236898
rect 573834 237454 574074 237486
rect 573834 237218 573836 237454
rect 574072 237218 574074 237454
rect 573834 237134 574074 237218
rect 573834 236898 573836 237134
rect 574072 236898 574074 237134
rect 573834 236866 574074 236898
rect 579288 237454 579888 237486
rect 579288 237218 579470 237454
rect 579706 237218 579888 237454
rect 579288 237134 579888 237218
rect 579288 236898 579470 237134
rect 579706 236898 579888 237134
rect 579288 236866 579888 236898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect 5200 219454 5800 219486
rect 5200 219218 5382 219454
rect 5618 219218 5800 219454
rect 5200 219134 5800 219218
rect 5200 218898 5382 219134
rect 5618 218898 5800 219134
rect 5200 218866 5800 218898
rect 12590 219454 12830 219486
rect 12590 219218 12592 219454
rect 12828 219218 12830 219454
rect 12590 219134 12830 219218
rect 12590 218898 12592 219134
rect 12828 218898 12830 219134
rect 12590 218866 12830 218898
rect 13436 219454 13676 219486
rect 13436 219218 13438 219454
rect 13674 219218 13676 219454
rect 13436 219134 13676 219218
rect 13436 218898 13438 219134
rect 13674 218898 13676 219134
rect 13436 218866 13676 218898
rect 22436 219454 22676 219486
rect 22436 219218 22438 219454
rect 22674 219218 22676 219454
rect 22436 219134 22676 219218
rect 22436 218898 22438 219134
rect 22674 218898 22676 219134
rect 22436 218866 22676 218898
rect 27226 219454 27466 219486
rect 27226 219218 27228 219454
rect 27464 219218 27466 219454
rect 27226 219134 27466 219218
rect 27226 218898 27228 219134
rect 27464 218898 27466 219134
rect 27226 218866 27466 218898
rect 28598 219454 28838 219486
rect 28598 219218 28600 219454
rect 28836 219218 28838 219454
rect 28598 219134 28838 219218
rect 28598 218898 28600 219134
rect 28836 218898 28838 219134
rect 28598 218866 28838 218898
rect 29444 219454 29684 219486
rect 29444 219218 29446 219454
rect 29682 219218 29684 219454
rect 29444 219134 29684 219218
rect 29444 218898 29446 219134
rect 29682 218898 29684 219134
rect 29444 218866 29684 218898
rect 38444 219454 38684 219486
rect 38444 219218 38446 219454
rect 38682 219218 38684 219454
rect 38444 219134 38684 219218
rect 38444 218898 38446 219134
rect 38682 218898 38684 219134
rect 38444 218866 38684 218898
rect 47444 219454 47684 219486
rect 47444 219218 47446 219454
rect 47682 219218 47684 219454
rect 47444 219134 47684 219218
rect 47444 218898 47446 219134
rect 47682 218898 47684 219134
rect 47444 218866 47684 218898
rect 56444 219454 56684 219486
rect 56444 219218 56446 219454
rect 56682 219218 56684 219454
rect 56444 219134 56684 219218
rect 56444 218898 56446 219134
rect 56682 218898 56684 219134
rect 56444 218866 56684 218898
rect 65444 219454 65684 219486
rect 65444 219218 65446 219454
rect 65682 219218 65684 219454
rect 65444 219134 65684 219218
rect 65444 218898 65446 219134
rect 65682 218898 65684 219134
rect 65444 218866 65684 218898
rect 67246 219454 67486 219486
rect 67246 219218 67248 219454
rect 67484 219218 67486 219454
rect 67246 219134 67486 219218
rect 67246 218898 67248 219134
rect 67484 218898 67486 219134
rect 67246 218866 67486 218898
rect 68618 219454 68858 219486
rect 68618 219218 68620 219454
rect 68856 219218 68858 219454
rect 68618 219134 68858 219218
rect 68618 218898 68620 219134
rect 68856 218898 68858 219134
rect 68618 218866 68858 218898
rect 69464 219454 69704 219486
rect 69464 219218 69466 219454
rect 69702 219218 69704 219454
rect 69464 219134 69704 219218
rect 69464 218898 69466 219134
rect 69702 218898 69704 219134
rect 69464 218866 69704 218898
rect 78464 219454 78704 219486
rect 78464 219218 78466 219454
rect 78702 219218 78704 219454
rect 78464 219134 78704 219218
rect 78464 218898 78466 219134
rect 78702 218898 78704 219134
rect 78464 218866 78704 218898
rect 87464 219454 87704 219486
rect 87464 219218 87466 219454
rect 87702 219218 87704 219454
rect 87464 219134 87704 219218
rect 87464 218898 87466 219134
rect 87702 218898 87704 219134
rect 87464 218866 87704 218898
rect 96464 219454 96704 219486
rect 96464 219218 96466 219454
rect 96702 219218 96704 219454
rect 96464 219134 96704 219218
rect 96464 218898 96466 219134
rect 96702 218898 96704 219134
rect 96464 218866 96704 218898
rect 105464 219454 105704 219486
rect 105464 219218 105466 219454
rect 105702 219218 105704 219454
rect 105464 219134 105704 219218
rect 105464 218898 105466 219134
rect 105702 218898 105704 219134
rect 105464 218866 105704 218898
rect 107266 219454 107506 219486
rect 107266 219218 107268 219454
rect 107504 219218 107506 219454
rect 107266 219134 107506 219218
rect 107266 218898 107268 219134
rect 107504 218898 107506 219134
rect 107266 218866 107506 218898
rect 108638 219454 108878 219486
rect 108638 219218 108640 219454
rect 108876 219218 108878 219454
rect 108638 219134 108878 219218
rect 108638 218898 108640 219134
rect 108876 218898 108878 219134
rect 108638 218866 108878 218898
rect 109484 219454 109724 219486
rect 109484 219218 109486 219454
rect 109722 219218 109724 219454
rect 109484 219134 109724 219218
rect 109484 218898 109486 219134
rect 109722 218898 109724 219134
rect 109484 218866 109724 218898
rect 118484 219454 118724 219486
rect 118484 219218 118486 219454
rect 118722 219218 118724 219454
rect 118484 219134 118724 219218
rect 118484 218898 118486 219134
rect 118722 218898 118724 219134
rect 118484 218866 118724 218898
rect 127484 219454 127724 219486
rect 127484 219218 127486 219454
rect 127722 219218 127724 219454
rect 127484 219134 127724 219218
rect 127484 218898 127486 219134
rect 127722 218898 127724 219134
rect 127484 218866 127724 218898
rect 136484 219454 136724 219486
rect 136484 219218 136486 219454
rect 136722 219218 136724 219454
rect 136484 219134 136724 219218
rect 136484 218898 136486 219134
rect 136722 218898 136724 219134
rect 136484 218866 136724 218898
rect 145484 219454 145724 219486
rect 145484 219218 145486 219454
rect 145722 219218 145724 219454
rect 145484 219134 145724 219218
rect 145484 218898 145486 219134
rect 145722 218898 145724 219134
rect 145484 218866 145724 218898
rect 147286 219454 147526 219486
rect 147286 219218 147288 219454
rect 147524 219218 147526 219454
rect 147286 219134 147526 219218
rect 147286 218898 147288 219134
rect 147524 218898 147526 219134
rect 147286 218866 147526 218898
rect 149658 219454 149898 219486
rect 149658 219218 149660 219454
rect 149896 219218 149898 219454
rect 149658 219134 149898 219218
rect 149658 218898 149660 219134
rect 149896 218898 149898 219134
rect 149658 218866 149898 218898
rect 150504 219454 150744 219486
rect 150504 219218 150506 219454
rect 150742 219218 150744 219454
rect 150504 219134 150744 219218
rect 150504 218898 150506 219134
rect 150742 218898 150744 219134
rect 150504 218866 150744 218898
rect 159504 219454 159744 219486
rect 159504 219218 159506 219454
rect 159742 219218 159744 219454
rect 159504 219134 159744 219218
rect 159504 218898 159506 219134
rect 159742 218898 159744 219134
rect 159504 218866 159744 218898
rect 168504 219454 168744 219486
rect 168504 219218 168506 219454
rect 168742 219218 168744 219454
rect 168504 219134 168744 219218
rect 168504 218898 168506 219134
rect 168742 218898 168744 219134
rect 168504 218866 168744 218898
rect 177504 219454 177744 219486
rect 177504 219218 177506 219454
rect 177742 219218 177744 219454
rect 177504 219134 177744 219218
rect 177504 218898 177506 219134
rect 177742 218898 177744 219134
rect 177504 218866 177744 218898
rect 186504 219454 186744 219486
rect 186504 219218 186506 219454
rect 186742 219218 186744 219454
rect 186504 219134 186744 219218
rect 186504 218898 186506 219134
rect 186742 218898 186744 219134
rect 186504 218866 186744 218898
rect 188306 219454 188546 219486
rect 188306 219218 188308 219454
rect 188544 219218 188546 219454
rect 188306 219134 188546 219218
rect 188306 218898 188308 219134
rect 188544 218898 188546 219134
rect 188306 218866 188546 218898
rect 190678 219454 190918 219486
rect 190678 219218 190680 219454
rect 190916 219218 190918 219454
rect 190678 219134 190918 219218
rect 190678 218898 190680 219134
rect 190916 218898 190918 219134
rect 190678 218866 190918 218898
rect 191524 219454 191764 219486
rect 191524 219218 191526 219454
rect 191762 219218 191764 219454
rect 191524 219134 191764 219218
rect 191524 218898 191526 219134
rect 191762 218898 191764 219134
rect 191524 218866 191764 218898
rect 200524 219454 200764 219486
rect 200524 219218 200526 219454
rect 200762 219218 200764 219454
rect 200524 219134 200764 219218
rect 200524 218898 200526 219134
rect 200762 218898 200764 219134
rect 200524 218866 200764 218898
rect 209524 219454 209764 219486
rect 209524 219218 209526 219454
rect 209762 219218 209764 219454
rect 209524 219134 209764 219218
rect 209524 218898 209526 219134
rect 209762 218898 209764 219134
rect 209524 218866 209764 218898
rect 218524 219454 218764 219486
rect 218524 219218 218526 219454
rect 218762 219218 218764 219454
rect 218524 219134 218764 219218
rect 218524 218898 218526 219134
rect 218762 218898 218764 219134
rect 218524 218866 218764 218898
rect 227524 219454 227764 219486
rect 227524 219218 227526 219454
rect 227762 219218 227764 219454
rect 227524 219134 227764 219218
rect 227524 218898 227526 219134
rect 227762 218898 227764 219134
rect 227524 218866 227764 218898
rect 229326 219454 229566 219486
rect 229326 219218 229328 219454
rect 229564 219218 229566 219454
rect 229326 219134 229566 219218
rect 229326 218898 229328 219134
rect 229564 218898 229566 219134
rect 229326 218866 229566 218898
rect 230698 219454 230938 219486
rect 230698 219218 230700 219454
rect 230936 219218 230938 219454
rect 230698 219134 230938 219218
rect 230698 218898 230700 219134
rect 230936 218898 230938 219134
rect 230698 218866 230938 218898
rect 231544 219454 231784 219486
rect 231544 219218 231546 219454
rect 231782 219218 231784 219454
rect 231544 219134 231784 219218
rect 231544 218898 231546 219134
rect 231782 218898 231784 219134
rect 231544 218866 231784 218898
rect 240544 219454 240784 219486
rect 240544 219218 240546 219454
rect 240782 219218 240784 219454
rect 240544 219134 240784 219218
rect 240544 218898 240546 219134
rect 240782 218898 240784 219134
rect 240544 218866 240784 218898
rect 249544 219454 249784 219486
rect 249544 219218 249546 219454
rect 249782 219218 249784 219454
rect 249544 219134 249784 219218
rect 249544 218898 249546 219134
rect 249782 218898 249784 219134
rect 249544 218866 249784 218898
rect 258544 219454 258784 219486
rect 258544 219218 258546 219454
rect 258782 219218 258784 219454
rect 258544 219134 258784 219218
rect 258544 218898 258546 219134
rect 258782 218898 258784 219134
rect 258544 218866 258784 218898
rect 267544 219454 267784 219486
rect 267544 219218 267546 219454
rect 267782 219218 267784 219454
rect 267544 219134 267784 219218
rect 267544 218898 267546 219134
rect 267782 218898 267784 219134
rect 267544 218866 267784 218898
rect 269346 219454 269586 219486
rect 269346 219218 269348 219454
rect 269584 219218 269586 219454
rect 269346 219134 269586 219218
rect 269346 218898 269348 219134
rect 269584 218898 269586 219134
rect 269346 218866 269586 218898
rect 270718 219454 270958 219486
rect 270718 219218 270720 219454
rect 270956 219218 270958 219454
rect 270718 219134 270958 219218
rect 270718 218898 270720 219134
rect 270956 218898 270958 219134
rect 270718 218866 270958 218898
rect 271564 219454 271804 219486
rect 271564 219218 271566 219454
rect 271802 219218 271804 219454
rect 271564 219134 271804 219218
rect 271564 218898 271566 219134
rect 271802 218898 271804 219134
rect 271564 218866 271804 218898
rect 280564 219454 280804 219486
rect 280564 219218 280566 219454
rect 280802 219218 280804 219454
rect 280564 219134 280804 219218
rect 280564 218898 280566 219134
rect 280802 218898 280804 219134
rect 280564 218866 280804 218898
rect 289564 219454 289804 219486
rect 289564 219218 289566 219454
rect 289802 219218 289804 219454
rect 289564 219134 289804 219218
rect 289564 218898 289566 219134
rect 289802 218898 289804 219134
rect 289564 218866 289804 218898
rect 298564 219454 298804 219486
rect 298564 219218 298566 219454
rect 298802 219218 298804 219454
rect 298564 219134 298804 219218
rect 298564 218898 298566 219134
rect 298802 218898 298804 219134
rect 298564 218866 298804 218898
rect 307564 219454 307804 219486
rect 307564 219218 307566 219454
rect 307802 219218 307804 219454
rect 307564 219134 307804 219218
rect 307564 218898 307566 219134
rect 307802 218898 307804 219134
rect 307564 218866 307804 218898
rect 309366 219454 309606 219486
rect 309366 219218 309368 219454
rect 309604 219218 309606 219454
rect 309366 219134 309606 219218
rect 309366 218898 309368 219134
rect 309604 218898 309606 219134
rect 309366 218866 309606 218898
rect 311738 219454 311978 219486
rect 311738 219218 311740 219454
rect 311976 219218 311978 219454
rect 311738 219134 311978 219218
rect 311738 218898 311740 219134
rect 311976 218898 311978 219134
rect 311738 218866 311978 218898
rect 312584 219454 312824 219486
rect 312584 219218 312586 219454
rect 312822 219218 312824 219454
rect 312584 219134 312824 219218
rect 312584 218898 312586 219134
rect 312822 218898 312824 219134
rect 312584 218866 312824 218898
rect 321584 219454 321824 219486
rect 321584 219218 321586 219454
rect 321822 219218 321824 219454
rect 321584 219134 321824 219218
rect 321584 218898 321586 219134
rect 321822 218898 321824 219134
rect 321584 218866 321824 218898
rect 330584 219454 330824 219486
rect 330584 219218 330586 219454
rect 330822 219218 330824 219454
rect 330584 219134 330824 219218
rect 330584 218898 330586 219134
rect 330822 218898 330824 219134
rect 330584 218866 330824 218898
rect 339584 219454 339824 219486
rect 339584 219218 339586 219454
rect 339822 219218 339824 219454
rect 339584 219134 339824 219218
rect 339584 218898 339586 219134
rect 339822 218898 339824 219134
rect 339584 218866 339824 218898
rect 348584 219454 348824 219486
rect 348584 219218 348586 219454
rect 348822 219218 348824 219454
rect 348584 219134 348824 219218
rect 348584 218898 348586 219134
rect 348822 218898 348824 219134
rect 348584 218866 348824 218898
rect 350386 219454 350626 219486
rect 350386 219218 350388 219454
rect 350624 219218 350626 219454
rect 350386 219134 350626 219218
rect 350386 218898 350388 219134
rect 350624 218898 350626 219134
rect 350386 218866 350626 218898
rect 352758 219454 352998 219486
rect 352758 219218 352760 219454
rect 352996 219218 352998 219454
rect 352758 219134 352998 219218
rect 352758 218898 352760 219134
rect 352996 218898 352998 219134
rect 352758 218866 352998 218898
rect 353604 219454 353844 219486
rect 353604 219218 353606 219454
rect 353842 219218 353844 219454
rect 353604 219134 353844 219218
rect 353604 218898 353606 219134
rect 353842 218898 353844 219134
rect 353604 218866 353844 218898
rect 362604 219454 362844 219486
rect 362604 219218 362606 219454
rect 362842 219218 362844 219454
rect 362604 219134 362844 219218
rect 362604 218898 362606 219134
rect 362842 218898 362844 219134
rect 362604 218866 362844 218898
rect 371604 219454 371844 219486
rect 371604 219218 371606 219454
rect 371842 219218 371844 219454
rect 371604 219134 371844 219218
rect 371604 218898 371606 219134
rect 371842 218898 371844 219134
rect 371604 218866 371844 218898
rect 380604 219454 380844 219486
rect 380604 219218 380606 219454
rect 380842 219218 380844 219454
rect 380604 219134 380844 219218
rect 380604 218898 380606 219134
rect 380842 218898 380844 219134
rect 380604 218866 380844 218898
rect 389604 219454 389844 219486
rect 389604 219218 389606 219454
rect 389842 219218 389844 219454
rect 389604 219134 389844 219218
rect 389604 218898 389606 219134
rect 389842 218898 389844 219134
rect 389604 218866 389844 218898
rect 391406 219454 391646 219486
rect 391406 219218 391408 219454
rect 391644 219218 391646 219454
rect 391406 219134 391646 219218
rect 391406 218898 391408 219134
rect 391644 218898 391646 219134
rect 391406 218866 391646 218898
rect 392778 219454 393018 219486
rect 392778 219218 392780 219454
rect 393016 219218 393018 219454
rect 392778 219134 393018 219218
rect 392778 218898 392780 219134
rect 393016 218898 393018 219134
rect 392778 218866 393018 218898
rect 393624 219454 393864 219486
rect 393624 219218 393626 219454
rect 393862 219218 393864 219454
rect 393624 219134 393864 219218
rect 393624 218898 393626 219134
rect 393862 218898 393864 219134
rect 393624 218866 393864 218898
rect 402624 219454 402864 219486
rect 402624 219218 402626 219454
rect 402862 219218 402864 219454
rect 402624 219134 402864 219218
rect 402624 218898 402626 219134
rect 402862 218898 402864 219134
rect 402624 218866 402864 218898
rect 411624 219454 411864 219486
rect 411624 219218 411626 219454
rect 411862 219218 411864 219454
rect 411624 219134 411864 219218
rect 411624 218898 411626 219134
rect 411862 218898 411864 219134
rect 411624 218866 411864 218898
rect 420624 219454 420864 219486
rect 420624 219218 420626 219454
rect 420862 219218 420864 219454
rect 420624 219134 420864 219218
rect 420624 218898 420626 219134
rect 420862 218898 420864 219134
rect 420624 218866 420864 218898
rect 429624 219454 429864 219486
rect 429624 219218 429626 219454
rect 429862 219218 429864 219454
rect 429624 219134 429864 219218
rect 429624 218898 429626 219134
rect 429862 218898 429864 219134
rect 429624 218866 429864 218898
rect 431426 219454 431666 219486
rect 431426 219218 431428 219454
rect 431664 219218 431666 219454
rect 431426 219134 431666 219218
rect 431426 218898 431428 219134
rect 431664 218898 431666 219134
rect 431426 218866 431666 218898
rect 432798 219454 433038 219486
rect 432798 219218 432800 219454
rect 433036 219218 433038 219454
rect 432798 219134 433038 219218
rect 432798 218898 432800 219134
rect 433036 218898 433038 219134
rect 432798 218866 433038 218898
rect 433644 219454 433884 219486
rect 433644 219218 433646 219454
rect 433882 219218 433884 219454
rect 433644 219134 433884 219218
rect 433644 218898 433646 219134
rect 433882 218898 433884 219134
rect 433644 218866 433884 218898
rect 442644 219454 442884 219486
rect 442644 219218 442646 219454
rect 442882 219218 442884 219454
rect 442644 219134 442884 219218
rect 442644 218898 442646 219134
rect 442882 218898 442884 219134
rect 442644 218866 442884 218898
rect 451644 219454 451884 219486
rect 451644 219218 451646 219454
rect 451882 219218 451884 219454
rect 451644 219134 451884 219218
rect 451644 218898 451646 219134
rect 451882 218898 451884 219134
rect 451644 218866 451884 218898
rect 460644 219454 460884 219486
rect 460644 219218 460646 219454
rect 460882 219218 460884 219454
rect 460644 219134 460884 219218
rect 460644 218898 460646 219134
rect 460882 218898 460884 219134
rect 460644 218866 460884 218898
rect 469644 219454 469884 219486
rect 469644 219218 469646 219454
rect 469882 219218 469884 219454
rect 469644 219134 469884 219218
rect 469644 218898 469646 219134
rect 469882 218898 469884 219134
rect 469644 218866 469884 218898
rect 471446 219454 471686 219486
rect 471446 219218 471448 219454
rect 471684 219218 471686 219454
rect 471446 219134 471686 219218
rect 471446 218898 471448 219134
rect 471684 218898 471686 219134
rect 471446 218866 471686 218898
rect 472818 219454 473058 219486
rect 472818 219218 472820 219454
rect 473056 219218 473058 219454
rect 472818 219134 473058 219218
rect 472818 218898 472820 219134
rect 473056 218898 473058 219134
rect 472818 218866 473058 218898
rect 473664 219454 473904 219486
rect 473664 219218 473666 219454
rect 473902 219218 473904 219454
rect 473664 219134 473904 219218
rect 473664 218898 473666 219134
rect 473902 218898 473904 219134
rect 473664 218866 473904 218898
rect 482664 219454 482904 219486
rect 482664 219218 482666 219454
rect 482902 219218 482904 219454
rect 482664 219134 482904 219218
rect 482664 218898 482666 219134
rect 482902 218898 482904 219134
rect 482664 218866 482904 218898
rect 491664 219454 491904 219486
rect 491664 219218 491666 219454
rect 491902 219218 491904 219454
rect 491664 219134 491904 219218
rect 491664 218898 491666 219134
rect 491902 218898 491904 219134
rect 491664 218866 491904 218898
rect 500664 219454 500904 219486
rect 500664 219218 500666 219454
rect 500902 219218 500904 219454
rect 500664 219134 500904 219218
rect 500664 218898 500666 219134
rect 500902 218898 500904 219134
rect 500664 218866 500904 218898
rect 509664 219454 509904 219486
rect 509664 219218 509666 219454
rect 509902 219218 509904 219454
rect 509664 219134 509904 219218
rect 509664 218898 509666 219134
rect 509902 218898 509904 219134
rect 509664 218866 509904 218898
rect 511466 219454 511706 219486
rect 511466 219218 511468 219454
rect 511704 219218 511706 219454
rect 511466 219134 511706 219218
rect 511466 218898 511468 219134
rect 511704 218898 511706 219134
rect 511466 218866 511706 218898
rect 512838 219454 513078 219486
rect 512838 219218 512840 219454
rect 513076 219218 513078 219454
rect 512838 219134 513078 219218
rect 512838 218898 512840 219134
rect 513076 218898 513078 219134
rect 512838 218866 513078 218898
rect 513684 219454 513924 219486
rect 513684 219218 513686 219454
rect 513922 219218 513924 219454
rect 513684 219134 513924 219218
rect 513684 218898 513686 219134
rect 513922 218898 513924 219134
rect 513684 218866 513924 218898
rect 522684 219454 522924 219486
rect 522684 219218 522686 219454
rect 522922 219218 522924 219454
rect 522684 219134 522924 219218
rect 522684 218898 522686 219134
rect 522922 218898 522924 219134
rect 522684 218866 522924 218898
rect 531684 219454 531924 219486
rect 531684 219218 531686 219454
rect 531922 219218 531924 219454
rect 531684 219134 531924 219218
rect 531684 218898 531686 219134
rect 531922 218898 531924 219134
rect 531684 218866 531924 218898
rect 540684 219454 540924 219486
rect 540684 219218 540686 219454
rect 540922 219218 540924 219454
rect 540684 219134 540924 219218
rect 540684 218898 540686 219134
rect 540922 218898 540924 219134
rect 540684 218866 540924 218898
rect 549684 219454 549924 219486
rect 549684 219218 549686 219454
rect 549922 219218 549924 219454
rect 549684 219134 549924 219218
rect 549684 218898 549686 219134
rect 549922 218898 549924 219134
rect 549684 218866 549924 218898
rect 551486 219454 551726 219486
rect 551486 219218 551488 219454
rect 551724 219218 551726 219454
rect 551486 219134 551726 219218
rect 551486 218898 551488 219134
rect 551724 218898 551726 219134
rect 551486 218866 551726 218898
rect 552858 219454 553098 219486
rect 552858 219218 552860 219454
rect 553096 219218 553098 219454
rect 552858 219134 553098 219218
rect 552858 218898 552860 219134
rect 553096 218898 553098 219134
rect 552858 218866 553098 218898
rect 553704 219454 553944 219486
rect 553704 219218 553706 219454
rect 553942 219218 553944 219454
rect 553704 219134 553944 219218
rect 553704 218898 553706 219134
rect 553942 218898 553944 219134
rect 553704 218866 553944 218898
rect 562704 219454 562944 219486
rect 562704 219218 562706 219454
rect 562942 219218 562944 219454
rect 562704 219134 562944 219218
rect 562704 218898 562706 219134
rect 562942 218898 562944 219134
rect 562704 218866 562944 218898
rect 571704 219454 571944 219486
rect 571704 219218 571706 219454
rect 571942 219218 571944 219454
rect 571704 219134 571944 219218
rect 571704 218898 571706 219134
rect 571942 218898 571944 219134
rect 571704 218866 571944 218898
rect 573474 219454 573714 219486
rect 573474 219218 573476 219454
rect 573712 219218 573714 219454
rect 573474 219134 573714 219218
rect 573474 218898 573476 219134
rect 573712 218898 573714 219134
rect 573474 218866 573714 218898
rect 578488 219454 579088 219486
rect 578488 219218 578670 219454
rect 578906 219218 579088 219454
rect 578488 219134 579088 219218
rect 578488 218898 578670 219134
rect 578906 218898 579088 219134
rect 578488 218866 579088 218898
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 4400 201454 5000 201486
rect 4400 201218 4582 201454
rect 4818 201218 5000 201454
rect 4400 201134 5000 201218
rect 4400 200898 4582 201134
rect 4818 200898 5000 201134
rect 4400 200866 5000 200898
rect 12230 201454 12470 201486
rect 12230 201218 12232 201454
rect 12468 201218 12470 201454
rect 12230 201134 12470 201218
rect 12230 200898 12232 201134
rect 12468 200898 12470 201134
rect 12230 200866 12470 200898
rect 13036 201454 13276 201486
rect 13036 201218 13038 201454
rect 13274 201218 13276 201454
rect 13036 201134 13276 201218
rect 13036 200898 13038 201134
rect 13274 200898 13276 201134
rect 13036 200866 13276 200898
rect 22036 201454 22276 201486
rect 22036 201218 22038 201454
rect 22274 201218 22276 201454
rect 22036 201134 22276 201218
rect 22036 200898 22038 201134
rect 22274 200898 22276 201134
rect 22036 200866 22276 200898
rect 27586 201454 27826 201486
rect 27586 201218 27588 201454
rect 27824 201218 27826 201454
rect 27586 201134 27826 201218
rect 27586 200898 27588 201134
rect 27824 200898 27826 201134
rect 27586 200866 27826 200898
rect 28238 201454 28478 201486
rect 28238 201218 28240 201454
rect 28476 201218 28478 201454
rect 28238 201134 28478 201218
rect 28238 200898 28240 201134
rect 28476 200898 28478 201134
rect 28238 200866 28478 200898
rect 29044 201454 29284 201486
rect 29044 201218 29046 201454
rect 29282 201218 29284 201454
rect 29044 201134 29284 201218
rect 29044 200898 29046 201134
rect 29282 200898 29284 201134
rect 29044 200866 29284 200898
rect 38044 201454 38284 201486
rect 38044 201218 38046 201454
rect 38282 201218 38284 201454
rect 38044 201134 38284 201218
rect 38044 200898 38046 201134
rect 38282 200898 38284 201134
rect 38044 200866 38284 200898
rect 47044 201454 47284 201486
rect 47044 201218 47046 201454
rect 47282 201218 47284 201454
rect 47044 201134 47284 201218
rect 47044 200898 47046 201134
rect 47282 200898 47284 201134
rect 47044 200866 47284 200898
rect 56044 201454 56284 201486
rect 56044 201218 56046 201454
rect 56282 201218 56284 201454
rect 56044 201134 56284 201218
rect 56044 200898 56046 201134
rect 56282 200898 56284 201134
rect 56044 200866 56284 200898
rect 65044 201454 65284 201486
rect 65044 201218 65046 201454
rect 65282 201218 65284 201454
rect 65044 201134 65284 201218
rect 65044 200898 65046 201134
rect 65282 200898 65284 201134
rect 65044 200866 65284 200898
rect 67606 201454 67846 201486
rect 67606 201218 67608 201454
rect 67844 201218 67846 201454
rect 67606 201134 67846 201218
rect 67606 200898 67608 201134
rect 67844 200898 67846 201134
rect 67606 200866 67846 200898
rect 68258 201454 68498 201486
rect 68258 201218 68260 201454
rect 68496 201218 68498 201454
rect 68258 201134 68498 201218
rect 68258 200898 68260 201134
rect 68496 200898 68498 201134
rect 68258 200866 68498 200898
rect 69064 201454 69304 201486
rect 69064 201218 69066 201454
rect 69302 201218 69304 201454
rect 69064 201134 69304 201218
rect 69064 200898 69066 201134
rect 69302 200898 69304 201134
rect 69064 200866 69304 200898
rect 78064 201454 78304 201486
rect 78064 201218 78066 201454
rect 78302 201218 78304 201454
rect 78064 201134 78304 201218
rect 78064 200898 78066 201134
rect 78302 200898 78304 201134
rect 78064 200866 78304 200898
rect 87064 201454 87304 201486
rect 87064 201218 87066 201454
rect 87302 201218 87304 201454
rect 87064 201134 87304 201218
rect 87064 200898 87066 201134
rect 87302 200898 87304 201134
rect 87064 200866 87304 200898
rect 96064 201454 96304 201486
rect 96064 201218 96066 201454
rect 96302 201218 96304 201454
rect 96064 201134 96304 201218
rect 96064 200898 96066 201134
rect 96302 200898 96304 201134
rect 96064 200866 96304 200898
rect 105064 201454 105304 201486
rect 105064 201218 105066 201454
rect 105302 201218 105304 201454
rect 105064 201134 105304 201218
rect 105064 200898 105066 201134
rect 105302 200898 105304 201134
rect 105064 200866 105304 200898
rect 107626 201454 107866 201486
rect 107626 201218 107628 201454
rect 107864 201218 107866 201454
rect 107626 201134 107866 201218
rect 107626 200898 107628 201134
rect 107864 200898 107866 201134
rect 107626 200866 107866 200898
rect 108278 201454 108518 201486
rect 108278 201218 108280 201454
rect 108516 201218 108518 201454
rect 108278 201134 108518 201218
rect 108278 200898 108280 201134
rect 108516 200898 108518 201134
rect 108278 200866 108518 200898
rect 109084 201454 109324 201486
rect 109084 201218 109086 201454
rect 109322 201218 109324 201454
rect 109084 201134 109324 201218
rect 109084 200898 109086 201134
rect 109322 200898 109324 201134
rect 109084 200866 109324 200898
rect 118084 201454 118324 201486
rect 118084 201218 118086 201454
rect 118322 201218 118324 201454
rect 118084 201134 118324 201218
rect 118084 200898 118086 201134
rect 118322 200898 118324 201134
rect 118084 200866 118324 200898
rect 127084 201454 127324 201486
rect 127084 201218 127086 201454
rect 127322 201218 127324 201454
rect 127084 201134 127324 201218
rect 127084 200898 127086 201134
rect 127322 200898 127324 201134
rect 127084 200866 127324 200898
rect 136084 201454 136324 201486
rect 136084 201218 136086 201454
rect 136322 201218 136324 201454
rect 136084 201134 136324 201218
rect 136084 200898 136086 201134
rect 136322 200898 136324 201134
rect 136084 200866 136324 200898
rect 145084 201454 145324 201486
rect 145084 201218 145086 201454
rect 145322 201218 145324 201454
rect 145084 201134 145324 201218
rect 145084 200898 145086 201134
rect 145322 200898 145324 201134
rect 145084 200866 145324 200898
rect 147646 201454 147886 201486
rect 147646 201218 147648 201454
rect 147884 201218 147886 201454
rect 147646 201134 147886 201218
rect 147646 200898 147648 201134
rect 147884 200898 147886 201134
rect 147646 200866 147886 200898
rect 149298 201454 149538 201486
rect 149298 201218 149300 201454
rect 149536 201218 149538 201454
rect 149298 201134 149538 201218
rect 149298 200898 149300 201134
rect 149536 200898 149538 201134
rect 149298 200866 149538 200898
rect 150104 201454 150344 201486
rect 150104 201218 150106 201454
rect 150342 201218 150344 201454
rect 150104 201134 150344 201218
rect 150104 200898 150106 201134
rect 150342 200898 150344 201134
rect 150104 200866 150344 200898
rect 159104 201454 159344 201486
rect 159104 201218 159106 201454
rect 159342 201218 159344 201454
rect 159104 201134 159344 201218
rect 159104 200898 159106 201134
rect 159342 200898 159344 201134
rect 159104 200866 159344 200898
rect 168104 201454 168344 201486
rect 168104 201218 168106 201454
rect 168342 201218 168344 201454
rect 168104 201134 168344 201218
rect 168104 200898 168106 201134
rect 168342 200898 168344 201134
rect 168104 200866 168344 200898
rect 177104 201454 177344 201486
rect 177104 201218 177106 201454
rect 177342 201218 177344 201454
rect 177104 201134 177344 201218
rect 177104 200898 177106 201134
rect 177342 200898 177344 201134
rect 177104 200866 177344 200898
rect 186104 201454 186344 201486
rect 186104 201218 186106 201454
rect 186342 201218 186344 201454
rect 186104 201134 186344 201218
rect 186104 200898 186106 201134
rect 186342 200898 186344 201134
rect 186104 200866 186344 200898
rect 188666 201454 188906 201486
rect 188666 201218 188668 201454
rect 188904 201218 188906 201454
rect 188666 201134 188906 201218
rect 188666 200898 188668 201134
rect 188904 200898 188906 201134
rect 188666 200866 188906 200898
rect 190318 201454 190558 201486
rect 190318 201218 190320 201454
rect 190556 201218 190558 201454
rect 190318 201134 190558 201218
rect 190318 200898 190320 201134
rect 190556 200898 190558 201134
rect 190318 200866 190558 200898
rect 191124 201454 191364 201486
rect 191124 201218 191126 201454
rect 191362 201218 191364 201454
rect 191124 201134 191364 201218
rect 191124 200898 191126 201134
rect 191362 200898 191364 201134
rect 191124 200866 191364 200898
rect 200124 201454 200364 201486
rect 200124 201218 200126 201454
rect 200362 201218 200364 201454
rect 200124 201134 200364 201218
rect 200124 200898 200126 201134
rect 200362 200898 200364 201134
rect 200124 200866 200364 200898
rect 209124 201454 209364 201486
rect 209124 201218 209126 201454
rect 209362 201218 209364 201454
rect 209124 201134 209364 201218
rect 209124 200898 209126 201134
rect 209362 200898 209364 201134
rect 209124 200866 209364 200898
rect 218124 201454 218364 201486
rect 218124 201218 218126 201454
rect 218362 201218 218364 201454
rect 218124 201134 218364 201218
rect 218124 200898 218126 201134
rect 218362 200898 218364 201134
rect 218124 200866 218364 200898
rect 227124 201454 227364 201486
rect 227124 201218 227126 201454
rect 227362 201218 227364 201454
rect 227124 201134 227364 201218
rect 227124 200898 227126 201134
rect 227362 200898 227364 201134
rect 227124 200866 227364 200898
rect 229686 201454 229926 201486
rect 229686 201218 229688 201454
rect 229924 201218 229926 201454
rect 229686 201134 229926 201218
rect 229686 200898 229688 201134
rect 229924 200898 229926 201134
rect 229686 200866 229926 200898
rect 230338 201454 230578 201486
rect 230338 201218 230340 201454
rect 230576 201218 230578 201454
rect 230338 201134 230578 201218
rect 230338 200898 230340 201134
rect 230576 200898 230578 201134
rect 230338 200866 230578 200898
rect 231144 201454 231384 201486
rect 231144 201218 231146 201454
rect 231382 201218 231384 201454
rect 231144 201134 231384 201218
rect 231144 200898 231146 201134
rect 231382 200898 231384 201134
rect 231144 200866 231384 200898
rect 240144 201454 240384 201486
rect 240144 201218 240146 201454
rect 240382 201218 240384 201454
rect 240144 201134 240384 201218
rect 240144 200898 240146 201134
rect 240382 200898 240384 201134
rect 240144 200866 240384 200898
rect 249144 201454 249384 201486
rect 249144 201218 249146 201454
rect 249382 201218 249384 201454
rect 249144 201134 249384 201218
rect 249144 200898 249146 201134
rect 249382 200898 249384 201134
rect 249144 200866 249384 200898
rect 258144 201454 258384 201486
rect 258144 201218 258146 201454
rect 258382 201218 258384 201454
rect 258144 201134 258384 201218
rect 258144 200898 258146 201134
rect 258382 200898 258384 201134
rect 258144 200866 258384 200898
rect 267144 201454 267384 201486
rect 267144 201218 267146 201454
rect 267382 201218 267384 201454
rect 267144 201134 267384 201218
rect 267144 200898 267146 201134
rect 267382 200898 267384 201134
rect 267144 200866 267384 200898
rect 269706 201454 269946 201486
rect 269706 201218 269708 201454
rect 269944 201218 269946 201454
rect 269706 201134 269946 201218
rect 269706 200898 269708 201134
rect 269944 200898 269946 201134
rect 269706 200866 269946 200898
rect 270358 201454 270598 201486
rect 270358 201218 270360 201454
rect 270596 201218 270598 201454
rect 270358 201134 270598 201218
rect 270358 200898 270360 201134
rect 270596 200898 270598 201134
rect 270358 200866 270598 200898
rect 271164 201454 271404 201486
rect 271164 201218 271166 201454
rect 271402 201218 271404 201454
rect 271164 201134 271404 201218
rect 271164 200898 271166 201134
rect 271402 200898 271404 201134
rect 271164 200866 271404 200898
rect 280164 201454 280404 201486
rect 280164 201218 280166 201454
rect 280402 201218 280404 201454
rect 280164 201134 280404 201218
rect 280164 200898 280166 201134
rect 280402 200898 280404 201134
rect 280164 200866 280404 200898
rect 289164 201454 289404 201486
rect 289164 201218 289166 201454
rect 289402 201218 289404 201454
rect 289164 201134 289404 201218
rect 289164 200898 289166 201134
rect 289402 200898 289404 201134
rect 289164 200866 289404 200898
rect 298164 201454 298404 201486
rect 298164 201218 298166 201454
rect 298402 201218 298404 201454
rect 298164 201134 298404 201218
rect 298164 200898 298166 201134
rect 298402 200898 298404 201134
rect 298164 200866 298404 200898
rect 307164 201454 307404 201486
rect 307164 201218 307166 201454
rect 307402 201218 307404 201454
rect 307164 201134 307404 201218
rect 307164 200898 307166 201134
rect 307402 200898 307404 201134
rect 307164 200866 307404 200898
rect 309726 201454 309966 201486
rect 309726 201218 309728 201454
rect 309964 201218 309966 201454
rect 309726 201134 309966 201218
rect 309726 200898 309728 201134
rect 309964 200898 309966 201134
rect 309726 200866 309966 200898
rect 311378 201454 311618 201486
rect 311378 201218 311380 201454
rect 311616 201218 311618 201454
rect 311378 201134 311618 201218
rect 311378 200898 311380 201134
rect 311616 200898 311618 201134
rect 311378 200866 311618 200898
rect 312184 201454 312424 201486
rect 312184 201218 312186 201454
rect 312422 201218 312424 201454
rect 312184 201134 312424 201218
rect 312184 200898 312186 201134
rect 312422 200898 312424 201134
rect 312184 200866 312424 200898
rect 321184 201454 321424 201486
rect 321184 201218 321186 201454
rect 321422 201218 321424 201454
rect 321184 201134 321424 201218
rect 321184 200898 321186 201134
rect 321422 200898 321424 201134
rect 321184 200866 321424 200898
rect 330184 201454 330424 201486
rect 330184 201218 330186 201454
rect 330422 201218 330424 201454
rect 330184 201134 330424 201218
rect 330184 200898 330186 201134
rect 330422 200898 330424 201134
rect 330184 200866 330424 200898
rect 339184 201454 339424 201486
rect 339184 201218 339186 201454
rect 339422 201218 339424 201454
rect 339184 201134 339424 201218
rect 339184 200898 339186 201134
rect 339422 200898 339424 201134
rect 339184 200866 339424 200898
rect 348184 201454 348424 201486
rect 348184 201218 348186 201454
rect 348422 201218 348424 201454
rect 348184 201134 348424 201218
rect 348184 200898 348186 201134
rect 348422 200898 348424 201134
rect 348184 200866 348424 200898
rect 350746 201454 350986 201486
rect 350746 201218 350748 201454
rect 350984 201218 350986 201454
rect 350746 201134 350986 201218
rect 350746 200898 350748 201134
rect 350984 200898 350986 201134
rect 350746 200866 350986 200898
rect 352398 201454 352638 201486
rect 352398 201218 352400 201454
rect 352636 201218 352638 201454
rect 352398 201134 352638 201218
rect 352398 200898 352400 201134
rect 352636 200898 352638 201134
rect 352398 200866 352638 200898
rect 353204 201454 353444 201486
rect 353204 201218 353206 201454
rect 353442 201218 353444 201454
rect 353204 201134 353444 201218
rect 353204 200898 353206 201134
rect 353442 200898 353444 201134
rect 353204 200866 353444 200898
rect 362204 201454 362444 201486
rect 362204 201218 362206 201454
rect 362442 201218 362444 201454
rect 362204 201134 362444 201218
rect 362204 200898 362206 201134
rect 362442 200898 362444 201134
rect 362204 200866 362444 200898
rect 371204 201454 371444 201486
rect 371204 201218 371206 201454
rect 371442 201218 371444 201454
rect 371204 201134 371444 201218
rect 371204 200898 371206 201134
rect 371442 200898 371444 201134
rect 371204 200866 371444 200898
rect 380204 201454 380444 201486
rect 380204 201218 380206 201454
rect 380442 201218 380444 201454
rect 380204 201134 380444 201218
rect 380204 200898 380206 201134
rect 380442 200898 380444 201134
rect 380204 200866 380444 200898
rect 389204 201454 389444 201486
rect 389204 201218 389206 201454
rect 389442 201218 389444 201454
rect 389204 201134 389444 201218
rect 389204 200898 389206 201134
rect 389442 200898 389444 201134
rect 389204 200866 389444 200898
rect 391766 201454 392006 201486
rect 391766 201218 391768 201454
rect 392004 201218 392006 201454
rect 391766 201134 392006 201218
rect 391766 200898 391768 201134
rect 392004 200898 392006 201134
rect 391766 200866 392006 200898
rect 392418 201454 392658 201486
rect 392418 201218 392420 201454
rect 392656 201218 392658 201454
rect 392418 201134 392658 201218
rect 392418 200898 392420 201134
rect 392656 200898 392658 201134
rect 392418 200866 392658 200898
rect 393224 201454 393464 201486
rect 393224 201218 393226 201454
rect 393462 201218 393464 201454
rect 393224 201134 393464 201218
rect 393224 200898 393226 201134
rect 393462 200898 393464 201134
rect 393224 200866 393464 200898
rect 402224 201454 402464 201486
rect 402224 201218 402226 201454
rect 402462 201218 402464 201454
rect 402224 201134 402464 201218
rect 402224 200898 402226 201134
rect 402462 200898 402464 201134
rect 402224 200866 402464 200898
rect 411224 201454 411464 201486
rect 411224 201218 411226 201454
rect 411462 201218 411464 201454
rect 411224 201134 411464 201218
rect 411224 200898 411226 201134
rect 411462 200898 411464 201134
rect 411224 200866 411464 200898
rect 420224 201454 420464 201486
rect 420224 201218 420226 201454
rect 420462 201218 420464 201454
rect 420224 201134 420464 201218
rect 420224 200898 420226 201134
rect 420462 200898 420464 201134
rect 420224 200866 420464 200898
rect 429224 201454 429464 201486
rect 429224 201218 429226 201454
rect 429462 201218 429464 201454
rect 429224 201134 429464 201218
rect 429224 200898 429226 201134
rect 429462 200898 429464 201134
rect 429224 200866 429464 200898
rect 431786 201454 432026 201486
rect 431786 201218 431788 201454
rect 432024 201218 432026 201454
rect 431786 201134 432026 201218
rect 431786 200898 431788 201134
rect 432024 200898 432026 201134
rect 431786 200866 432026 200898
rect 432438 201454 432678 201486
rect 432438 201218 432440 201454
rect 432676 201218 432678 201454
rect 432438 201134 432678 201218
rect 432438 200898 432440 201134
rect 432676 200898 432678 201134
rect 432438 200866 432678 200898
rect 433244 201454 433484 201486
rect 433244 201218 433246 201454
rect 433482 201218 433484 201454
rect 433244 201134 433484 201218
rect 433244 200898 433246 201134
rect 433482 200898 433484 201134
rect 433244 200866 433484 200898
rect 442244 201454 442484 201486
rect 442244 201218 442246 201454
rect 442482 201218 442484 201454
rect 442244 201134 442484 201218
rect 442244 200898 442246 201134
rect 442482 200898 442484 201134
rect 442244 200866 442484 200898
rect 451244 201454 451484 201486
rect 451244 201218 451246 201454
rect 451482 201218 451484 201454
rect 451244 201134 451484 201218
rect 451244 200898 451246 201134
rect 451482 200898 451484 201134
rect 451244 200866 451484 200898
rect 460244 201454 460484 201486
rect 460244 201218 460246 201454
rect 460482 201218 460484 201454
rect 460244 201134 460484 201218
rect 460244 200898 460246 201134
rect 460482 200898 460484 201134
rect 460244 200866 460484 200898
rect 469244 201454 469484 201486
rect 469244 201218 469246 201454
rect 469482 201218 469484 201454
rect 469244 201134 469484 201218
rect 469244 200898 469246 201134
rect 469482 200898 469484 201134
rect 469244 200866 469484 200898
rect 471806 201454 472046 201486
rect 471806 201218 471808 201454
rect 472044 201218 472046 201454
rect 471806 201134 472046 201218
rect 471806 200898 471808 201134
rect 472044 200898 472046 201134
rect 471806 200866 472046 200898
rect 472458 201454 472698 201486
rect 472458 201218 472460 201454
rect 472696 201218 472698 201454
rect 472458 201134 472698 201218
rect 472458 200898 472460 201134
rect 472696 200898 472698 201134
rect 472458 200866 472698 200898
rect 473264 201454 473504 201486
rect 473264 201218 473266 201454
rect 473502 201218 473504 201454
rect 473264 201134 473504 201218
rect 473264 200898 473266 201134
rect 473502 200898 473504 201134
rect 473264 200866 473504 200898
rect 482264 201454 482504 201486
rect 482264 201218 482266 201454
rect 482502 201218 482504 201454
rect 482264 201134 482504 201218
rect 482264 200898 482266 201134
rect 482502 200898 482504 201134
rect 482264 200866 482504 200898
rect 491264 201454 491504 201486
rect 491264 201218 491266 201454
rect 491502 201218 491504 201454
rect 491264 201134 491504 201218
rect 491264 200898 491266 201134
rect 491502 200898 491504 201134
rect 491264 200866 491504 200898
rect 500264 201454 500504 201486
rect 500264 201218 500266 201454
rect 500502 201218 500504 201454
rect 500264 201134 500504 201218
rect 500264 200898 500266 201134
rect 500502 200898 500504 201134
rect 500264 200866 500504 200898
rect 509264 201454 509504 201486
rect 509264 201218 509266 201454
rect 509502 201218 509504 201454
rect 509264 201134 509504 201218
rect 509264 200898 509266 201134
rect 509502 200898 509504 201134
rect 509264 200866 509504 200898
rect 511826 201454 512066 201486
rect 511826 201218 511828 201454
rect 512064 201218 512066 201454
rect 511826 201134 512066 201218
rect 511826 200898 511828 201134
rect 512064 200898 512066 201134
rect 511826 200866 512066 200898
rect 512478 201454 512718 201486
rect 512478 201218 512480 201454
rect 512716 201218 512718 201454
rect 512478 201134 512718 201218
rect 512478 200898 512480 201134
rect 512716 200898 512718 201134
rect 512478 200866 512718 200898
rect 513284 201454 513524 201486
rect 513284 201218 513286 201454
rect 513522 201218 513524 201454
rect 513284 201134 513524 201218
rect 513284 200898 513286 201134
rect 513522 200898 513524 201134
rect 513284 200866 513524 200898
rect 522284 201454 522524 201486
rect 522284 201218 522286 201454
rect 522522 201218 522524 201454
rect 522284 201134 522524 201218
rect 522284 200898 522286 201134
rect 522522 200898 522524 201134
rect 522284 200866 522524 200898
rect 531284 201454 531524 201486
rect 531284 201218 531286 201454
rect 531522 201218 531524 201454
rect 531284 201134 531524 201218
rect 531284 200898 531286 201134
rect 531522 200898 531524 201134
rect 531284 200866 531524 200898
rect 540284 201454 540524 201486
rect 540284 201218 540286 201454
rect 540522 201218 540524 201454
rect 540284 201134 540524 201218
rect 540284 200898 540286 201134
rect 540522 200898 540524 201134
rect 540284 200866 540524 200898
rect 549284 201454 549524 201486
rect 549284 201218 549286 201454
rect 549522 201218 549524 201454
rect 549284 201134 549524 201218
rect 549284 200898 549286 201134
rect 549522 200898 549524 201134
rect 549284 200866 549524 200898
rect 551846 201454 552086 201486
rect 551846 201218 551848 201454
rect 552084 201218 552086 201454
rect 551846 201134 552086 201218
rect 551846 200898 551848 201134
rect 552084 200898 552086 201134
rect 551846 200866 552086 200898
rect 552498 201454 552738 201486
rect 552498 201218 552500 201454
rect 552736 201218 552738 201454
rect 552498 201134 552738 201218
rect 552498 200898 552500 201134
rect 552736 200898 552738 201134
rect 552498 200866 552738 200898
rect 553304 201454 553544 201486
rect 553304 201218 553306 201454
rect 553542 201218 553544 201454
rect 553304 201134 553544 201218
rect 553304 200898 553306 201134
rect 553542 200898 553544 201134
rect 553304 200866 553544 200898
rect 562304 201454 562544 201486
rect 562304 201218 562306 201454
rect 562542 201218 562544 201454
rect 562304 201134 562544 201218
rect 562304 200898 562306 201134
rect 562542 200898 562544 201134
rect 562304 200866 562544 200898
rect 571304 201454 571544 201486
rect 571304 201218 571306 201454
rect 571542 201218 571544 201454
rect 571304 201134 571544 201218
rect 571304 200898 571306 201134
rect 571542 200898 571544 201134
rect 571304 200866 571544 200898
rect 573834 201454 574074 201486
rect 573834 201218 573836 201454
rect 574072 201218 574074 201454
rect 573834 201134 574074 201218
rect 573834 200898 573836 201134
rect 574072 200898 574074 201134
rect 573834 200866 574074 200898
rect 579288 201454 579888 201486
rect 579288 201218 579470 201454
rect 579706 201218 579888 201454
rect 579288 201134 579888 201218
rect 579288 200898 579470 201134
rect 579706 200898 579888 201134
rect 579288 200866 579888 200898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect 5200 183454 5800 183486
rect 5200 183218 5382 183454
rect 5618 183218 5800 183454
rect 5200 183134 5800 183218
rect 5200 182898 5382 183134
rect 5618 182898 5800 183134
rect 5200 182866 5800 182898
rect 12590 183454 12830 183486
rect 12590 183218 12592 183454
rect 12828 183218 12830 183454
rect 12590 183134 12830 183218
rect 12590 182898 12592 183134
rect 12828 182898 12830 183134
rect 12590 182866 12830 182898
rect 13436 183454 13676 183486
rect 13436 183218 13438 183454
rect 13674 183218 13676 183454
rect 13436 183134 13676 183218
rect 13436 182898 13438 183134
rect 13674 182898 13676 183134
rect 13436 182866 13676 182898
rect 22436 183454 22676 183486
rect 22436 183218 22438 183454
rect 22674 183218 22676 183454
rect 22436 183134 22676 183218
rect 22436 182898 22438 183134
rect 22674 182898 22676 183134
rect 22436 182866 22676 182898
rect 27226 183454 27466 183486
rect 27226 183218 27228 183454
rect 27464 183218 27466 183454
rect 27226 183134 27466 183218
rect 27226 182898 27228 183134
rect 27464 182898 27466 183134
rect 27226 182866 27466 182898
rect 28598 183454 28838 183486
rect 28598 183218 28600 183454
rect 28836 183218 28838 183454
rect 28598 183134 28838 183218
rect 28598 182898 28600 183134
rect 28836 182898 28838 183134
rect 28598 182866 28838 182898
rect 29444 183454 29684 183486
rect 29444 183218 29446 183454
rect 29682 183218 29684 183454
rect 29444 183134 29684 183218
rect 29444 182898 29446 183134
rect 29682 182898 29684 183134
rect 29444 182866 29684 182898
rect 38444 183454 38684 183486
rect 38444 183218 38446 183454
rect 38682 183218 38684 183454
rect 38444 183134 38684 183218
rect 38444 182898 38446 183134
rect 38682 182898 38684 183134
rect 38444 182866 38684 182898
rect 47444 183454 47684 183486
rect 47444 183218 47446 183454
rect 47682 183218 47684 183454
rect 47444 183134 47684 183218
rect 47444 182898 47446 183134
rect 47682 182898 47684 183134
rect 47444 182866 47684 182898
rect 56444 183454 56684 183486
rect 56444 183218 56446 183454
rect 56682 183218 56684 183454
rect 56444 183134 56684 183218
rect 56444 182898 56446 183134
rect 56682 182898 56684 183134
rect 56444 182866 56684 182898
rect 65444 183454 65684 183486
rect 65444 183218 65446 183454
rect 65682 183218 65684 183454
rect 65444 183134 65684 183218
rect 65444 182898 65446 183134
rect 65682 182898 65684 183134
rect 65444 182866 65684 182898
rect 67246 183454 67486 183486
rect 67246 183218 67248 183454
rect 67484 183218 67486 183454
rect 67246 183134 67486 183218
rect 67246 182898 67248 183134
rect 67484 182898 67486 183134
rect 67246 182866 67486 182898
rect 68618 183454 68858 183486
rect 68618 183218 68620 183454
rect 68856 183218 68858 183454
rect 68618 183134 68858 183218
rect 68618 182898 68620 183134
rect 68856 182898 68858 183134
rect 68618 182866 68858 182898
rect 69464 183454 69704 183486
rect 69464 183218 69466 183454
rect 69702 183218 69704 183454
rect 69464 183134 69704 183218
rect 69464 182898 69466 183134
rect 69702 182898 69704 183134
rect 69464 182866 69704 182898
rect 78464 183454 78704 183486
rect 78464 183218 78466 183454
rect 78702 183218 78704 183454
rect 78464 183134 78704 183218
rect 78464 182898 78466 183134
rect 78702 182898 78704 183134
rect 78464 182866 78704 182898
rect 87464 183454 87704 183486
rect 87464 183218 87466 183454
rect 87702 183218 87704 183454
rect 87464 183134 87704 183218
rect 87464 182898 87466 183134
rect 87702 182898 87704 183134
rect 87464 182866 87704 182898
rect 96464 183454 96704 183486
rect 96464 183218 96466 183454
rect 96702 183218 96704 183454
rect 96464 183134 96704 183218
rect 96464 182898 96466 183134
rect 96702 182898 96704 183134
rect 96464 182866 96704 182898
rect 105464 183454 105704 183486
rect 105464 183218 105466 183454
rect 105702 183218 105704 183454
rect 105464 183134 105704 183218
rect 105464 182898 105466 183134
rect 105702 182898 105704 183134
rect 105464 182866 105704 182898
rect 107266 183454 107506 183486
rect 107266 183218 107268 183454
rect 107504 183218 107506 183454
rect 107266 183134 107506 183218
rect 107266 182898 107268 183134
rect 107504 182898 107506 183134
rect 107266 182866 107506 182898
rect 108638 183454 108878 183486
rect 108638 183218 108640 183454
rect 108876 183218 108878 183454
rect 108638 183134 108878 183218
rect 108638 182898 108640 183134
rect 108876 182898 108878 183134
rect 108638 182866 108878 182898
rect 109484 183454 109724 183486
rect 109484 183218 109486 183454
rect 109722 183218 109724 183454
rect 109484 183134 109724 183218
rect 109484 182898 109486 183134
rect 109722 182898 109724 183134
rect 109484 182866 109724 182898
rect 118484 183454 118724 183486
rect 118484 183218 118486 183454
rect 118722 183218 118724 183454
rect 118484 183134 118724 183218
rect 118484 182898 118486 183134
rect 118722 182898 118724 183134
rect 118484 182866 118724 182898
rect 127484 183454 127724 183486
rect 127484 183218 127486 183454
rect 127722 183218 127724 183454
rect 127484 183134 127724 183218
rect 127484 182898 127486 183134
rect 127722 182898 127724 183134
rect 127484 182866 127724 182898
rect 136484 183454 136724 183486
rect 136484 183218 136486 183454
rect 136722 183218 136724 183454
rect 136484 183134 136724 183218
rect 136484 182898 136486 183134
rect 136722 182898 136724 183134
rect 136484 182866 136724 182898
rect 145484 183454 145724 183486
rect 145484 183218 145486 183454
rect 145722 183218 145724 183454
rect 145484 183134 145724 183218
rect 145484 182898 145486 183134
rect 145722 182898 145724 183134
rect 145484 182866 145724 182898
rect 147286 183454 147526 183486
rect 147286 183218 147288 183454
rect 147524 183218 147526 183454
rect 147286 183134 147526 183218
rect 147286 182898 147288 183134
rect 147524 182898 147526 183134
rect 147286 182866 147526 182898
rect 149658 183454 149898 183486
rect 149658 183218 149660 183454
rect 149896 183218 149898 183454
rect 149658 183134 149898 183218
rect 149658 182898 149660 183134
rect 149896 182898 149898 183134
rect 149658 182866 149898 182898
rect 150504 183454 150744 183486
rect 150504 183218 150506 183454
rect 150742 183218 150744 183454
rect 150504 183134 150744 183218
rect 150504 182898 150506 183134
rect 150742 182898 150744 183134
rect 150504 182866 150744 182898
rect 159504 183454 159744 183486
rect 159504 183218 159506 183454
rect 159742 183218 159744 183454
rect 159504 183134 159744 183218
rect 159504 182898 159506 183134
rect 159742 182898 159744 183134
rect 159504 182866 159744 182898
rect 168504 183454 168744 183486
rect 168504 183218 168506 183454
rect 168742 183218 168744 183454
rect 168504 183134 168744 183218
rect 168504 182898 168506 183134
rect 168742 182898 168744 183134
rect 168504 182866 168744 182898
rect 177504 183454 177744 183486
rect 177504 183218 177506 183454
rect 177742 183218 177744 183454
rect 177504 183134 177744 183218
rect 177504 182898 177506 183134
rect 177742 182898 177744 183134
rect 177504 182866 177744 182898
rect 186504 183454 186744 183486
rect 186504 183218 186506 183454
rect 186742 183218 186744 183454
rect 186504 183134 186744 183218
rect 186504 182898 186506 183134
rect 186742 182898 186744 183134
rect 186504 182866 186744 182898
rect 188306 183454 188546 183486
rect 188306 183218 188308 183454
rect 188544 183218 188546 183454
rect 188306 183134 188546 183218
rect 188306 182898 188308 183134
rect 188544 182898 188546 183134
rect 188306 182866 188546 182898
rect 190678 183454 190918 183486
rect 190678 183218 190680 183454
rect 190916 183218 190918 183454
rect 190678 183134 190918 183218
rect 190678 182898 190680 183134
rect 190916 182898 190918 183134
rect 190678 182866 190918 182898
rect 191524 183454 191764 183486
rect 191524 183218 191526 183454
rect 191762 183218 191764 183454
rect 191524 183134 191764 183218
rect 191524 182898 191526 183134
rect 191762 182898 191764 183134
rect 191524 182866 191764 182898
rect 200524 183454 200764 183486
rect 200524 183218 200526 183454
rect 200762 183218 200764 183454
rect 200524 183134 200764 183218
rect 200524 182898 200526 183134
rect 200762 182898 200764 183134
rect 200524 182866 200764 182898
rect 209524 183454 209764 183486
rect 209524 183218 209526 183454
rect 209762 183218 209764 183454
rect 209524 183134 209764 183218
rect 209524 182898 209526 183134
rect 209762 182898 209764 183134
rect 209524 182866 209764 182898
rect 218524 183454 218764 183486
rect 218524 183218 218526 183454
rect 218762 183218 218764 183454
rect 218524 183134 218764 183218
rect 218524 182898 218526 183134
rect 218762 182898 218764 183134
rect 218524 182866 218764 182898
rect 227524 183454 227764 183486
rect 227524 183218 227526 183454
rect 227762 183218 227764 183454
rect 227524 183134 227764 183218
rect 227524 182898 227526 183134
rect 227762 182898 227764 183134
rect 227524 182866 227764 182898
rect 229326 183454 229566 183486
rect 229326 183218 229328 183454
rect 229564 183218 229566 183454
rect 229326 183134 229566 183218
rect 229326 182898 229328 183134
rect 229564 182898 229566 183134
rect 229326 182866 229566 182898
rect 230698 183454 230938 183486
rect 230698 183218 230700 183454
rect 230936 183218 230938 183454
rect 230698 183134 230938 183218
rect 230698 182898 230700 183134
rect 230936 182898 230938 183134
rect 230698 182866 230938 182898
rect 231544 183454 231784 183486
rect 231544 183218 231546 183454
rect 231782 183218 231784 183454
rect 231544 183134 231784 183218
rect 231544 182898 231546 183134
rect 231782 182898 231784 183134
rect 231544 182866 231784 182898
rect 240544 183454 240784 183486
rect 240544 183218 240546 183454
rect 240782 183218 240784 183454
rect 240544 183134 240784 183218
rect 240544 182898 240546 183134
rect 240782 182898 240784 183134
rect 240544 182866 240784 182898
rect 249544 183454 249784 183486
rect 249544 183218 249546 183454
rect 249782 183218 249784 183454
rect 249544 183134 249784 183218
rect 249544 182898 249546 183134
rect 249782 182898 249784 183134
rect 249544 182866 249784 182898
rect 258544 183454 258784 183486
rect 258544 183218 258546 183454
rect 258782 183218 258784 183454
rect 258544 183134 258784 183218
rect 258544 182898 258546 183134
rect 258782 182898 258784 183134
rect 258544 182866 258784 182898
rect 267544 183454 267784 183486
rect 267544 183218 267546 183454
rect 267782 183218 267784 183454
rect 267544 183134 267784 183218
rect 267544 182898 267546 183134
rect 267782 182898 267784 183134
rect 267544 182866 267784 182898
rect 269346 183454 269586 183486
rect 269346 183218 269348 183454
rect 269584 183218 269586 183454
rect 269346 183134 269586 183218
rect 269346 182898 269348 183134
rect 269584 182898 269586 183134
rect 269346 182866 269586 182898
rect 270718 183454 270958 183486
rect 270718 183218 270720 183454
rect 270956 183218 270958 183454
rect 270718 183134 270958 183218
rect 270718 182898 270720 183134
rect 270956 182898 270958 183134
rect 270718 182866 270958 182898
rect 271564 183454 271804 183486
rect 271564 183218 271566 183454
rect 271802 183218 271804 183454
rect 271564 183134 271804 183218
rect 271564 182898 271566 183134
rect 271802 182898 271804 183134
rect 271564 182866 271804 182898
rect 280564 183454 280804 183486
rect 280564 183218 280566 183454
rect 280802 183218 280804 183454
rect 280564 183134 280804 183218
rect 280564 182898 280566 183134
rect 280802 182898 280804 183134
rect 280564 182866 280804 182898
rect 289564 183454 289804 183486
rect 289564 183218 289566 183454
rect 289802 183218 289804 183454
rect 289564 183134 289804 183218
rect 289564 182898 289566 183134
rect 289802 182898 289804 183134
rect 289564 182866 289804 182898
rect 298564 183454 298804 183486
rect 298564 183218 298566 183454
rect 298802 183218 298804 183454
rect 298564 183134 298804 183218
rect 298564 182898 298566 183134
rect 298802 182898 298804 183134
rect 298564 182866 298804 182898
rect 307564 183454 307804 183486
rect 307564 183218 307566 183454
rect 307802 183218 307804 183454
rect 307564 183134 307804 183218
rect 307564 182898 307566 183134
rect 307802 182898 307804 183134
rect 307564 182866 307804 182898
rect 309366 183454 309606 183486
rect 309366 183218 309368 183454
rect 309604 183218 309606 183454
rect 309366 183134 309606 183218
rect 309366 182898 309368 183134
rect 309604 182898 309606 183134
rect 309366 182866 309606 182898
rect 311738 183454 311978 183486
rect 311738 183218 311740 183454
rect 311976 183218 311978 183454
rect 311738 183134 311978 183218
rect 311738 182898 311740 183134
rect 311976 182898 311978 183134
rect 311738 182866 311978 182898
rect 312584 183454 312824 183486
rect 312584 183218 312586 183454
rect 312822 183218 312824 183454
rect 312584 183134 312824 183218
rect 312584 182898 312586 183134
rect 312822 182898 312824 183134
rect 312584 182866 312824 182898
rect 321584 183454 321824 183486
rect 321584 183218 321586 183454
rect 321822 183218 321824 183454
rect 321584 183134 321824 183218
rect 321584 182898 321586 183134
rect 321822 182898 321824 183134
rect 321584 182866 321824 182898
rect 330584 183454 330824 183486
rect 330584 183218 330586 183454
rect 330822 183218 330824 183454
rect 330584 183134 330824 183218
rect 330584 182898 330586 183134
rect 330822 182898 330824 183134
rect 330584 182866 330824 182898
rect 339584 183454 339824 183486
rect 339584 183218 339586 183454
rect 339822 183218 339824 183454
rect 339584 183134 339824 183218
rect 339584 182898 339586 183134
rect 339822 182898 339824 183134
rect 339584 182866 339824 182898
rect 348584 183454 348824 183486
rect 348584 183218 348586 183454
rect 348822 183218 348824 183454
rect 348584 183134 348824 183218
rect 348584 182898 348586 183134
rect 348822 182898 348824 183134
rect 348584 182866 348824 182898
rect 350386 183454 350626 183486
rect 350386 183218 350388 183454
rect 350624 183218 350626 183454
rect 350386 183134 350626 183218
rect 350386 182898 350388 183134
rect 350624 182898 350626 183134
rect 350386 182866 350626 182898
rect 352758 183454 352998 183486
rect 352758 183218 352760 183454
rect 352996 183218 352998 183454
rect 352758 183134 352998 183218
rect 352758 182898 352760 183134
rect 352996 182898 352998 183134
rect 352758 182866 352998 182898
rect 353604 183454 353844 183486
rect 353604 183218 353606 183454
rect 353842 183218 353844 183454
rect 353604 183134 353844 183218
rect 353604 182898 353606 183134
rect 353842 182898 353844 183134
rect 353604 182866 353844 182898
rect 362604 183454 362844 183486
rect 362604 183218 362606 183454
rect 362842 183218 362844 183454
rect 362604 183134 362844 183218
rect 362604 182898 362606 183134
rect 362842 182898 362844 183134
rect 362604 182866 362844 182898
rect 371604 183454 371844 183486
rect 371604 183218 371606 183454
rect 371842 183218 371844 183454
rect 371604 183134 371844 183218
rect 371604 182898 371606 183134
rect 371842 182898 371844 183134
rect 371604 182866 371844 182898
rect 380604 183454 380844 183486
rect 380604 183218 380606 183454
rect 380842 183218 380844 183454
rect 380604 183134 380844 183218
rect 380604 182898 380606 183134
rect 380842 182898 380844 183134
rect 380604 182866 380844 182898
rect 389604 183454 389844 183486
rect 389604 183218 389606 183454
rect 389842 183218 389844 183454
rect 389604 183134 389844 183218
rect 389604 182898 389606 183134
rect 389842 182898 389844 183134
rect 389604 182866 389844 182898
rect 391406 183454 391646 183486
rect 391406 183218 391408 183454
rect 391644 183218 391646 183454
rect 391406 183134 391646 183218
rect 391406 182898 391408 183134
rect 391644 182898 391646 183134
rect 391406 182866 391646 182898
rect 392778 183454 393018 183486
rect 392778 183218 392780 183454
rect 393016 183218 393018 183454
rect 392778 183134 393018 183218
rect 392778 182898 392780 183134
rect 393016 182898 393018 183134
rect 392778 182866 393018 182898
rect 393624 183454 393864 183486
rect 393624 183218 393626 183454
rect 393862 183218 393864 183454
rect 393624 183134 393864 183218
rect 393624 182898 393626 183134
rect 393862 182898 393864 183134
rect 393624 182866 393864 182898
rect 402624 183454 402864 183486
rect 402624 183218 402626 183454
rect 402862 183218 402864 183454
rect 402624 183134 402864 183218
rect 402624 182898 402626 183134
rect 402862 182898 402864 183134
rect 402624 182866 402864 182898
rect 411624 183454 411864 183486
rect 411624 183218 411626 183454
rect 411862 183218 411864 183454
rect 411624 183134 411864 183218
rect 411624 182898 411626 183134
rect 411862 182898 411864 183134
rect 411624 182866 411864 182898
rect 420624 183454 420864 183486
rect 420624 183218 420626 183454
rect 420862 183218 420864 183454
rect 420624 183134 420864 183218
rect 420624 182898 420626 183134
rect 420862 182898 420864 183134
rect 420624 182866 420864 182898
rect 429624 183454 429864 183486
rect 429624 183218 429626 183454
rect 429862 183218 429864 183454
rect 429624 183134 429864 183218
rect 429624 182898 429626 183134
rect 429862 182898 429864 183134
rect 429624 182866 429864 182898
rect 431426 183454 431666 183486
rect 431426 183218 431428 183454
rect 431664 183218 431666 183454
rect 431426 183134 431666 183218
rect 431426 182898 431428 183134
rect 431664 182898 431666 183134
rect 431426 182866 431666 182898
rect 432798 183454 433038 183486
rect 432798 183218 432800 183454
rect 433036 183218 433038 183454
rect 432798 183134 433038 183218
rect 432798 182898 432800 183134
rect 433036 182898 433038 183134
rect 432798 182866 433038 182898
rect 433644 183454 433884 183486
rect 433644 183218 433646 183454
rect 433882 183218 433884 183454
rect 433644 183134 433884 183218
rect 433644 182898 433646 183134
rect 433882 182898 433884 183134
rect 433644 182866 433884 182898
rect 442644 183454 442884 183486
rect 442644 183218 442646 183454
rect 442882 183218 442884 183454
rect 442644 183134 442884 183218
rect 442644 182898 442646 183134
rect 442882 182898 442884 183134
rect 442644 182866 442884 182898
rect 451644 183454 451884 183486
rect 451644 183218 451646 183454
rect 451882 183218 451884 183454
rect 451644 183134 451884 183218
rect 451644 182898 451646 183134
rect 451882 182898 451884 183134
rect 451644 182866 451884 182898
rect 460644 183454 460884 183486
rect 460644 183218 460646 183454
rect 460882 183218 460884 183454
rect 460644 183134 460884 183218
rect 460644 182898 460646 183134
rect 460882 182898 460884 183134
rect 460644 182866 460884 182898
rect 469644 183454 469884 183486
rect 469644 183218 469646 183454
rect 469882 183218 469884 183454
rect 469644 183134 469884 183218
rect 469644 182898 469646 183134
rect 469882 182898 469884 183134
rect 469644 182866 469884 182898
rect 471446 183454 471686 183486
rect 471446 183218 471448 183454
rect 471684 183218 471686 183454
rect 471446 183134 471686 183218
rect 471446 182898 471448 183134
rect 471684 182898 471686 183134
rect 471446 182866 471686 182898
rect 472818 183454 473058 183486
rect 472818 183218 472820 183454
rect 473056 183218 473058 183454
rect 472818 183134 473058 183218
rect 472818 182898 472820 183134
rect 473056 182898 473058 183134
rect 472818 182866 473058 182898
rect 473664 183454 473904 183486
rect 473664 183218 473666 183454
rect 473902 183218 473904 183454
rect 473664 183134 473904 183218
rect 473664 182898 473666 183134
rect 473902 182898 473904 183134
rect 473664 182866 473904 182898
rect 482664 183454 482904 183486
rect 482664 183218 482666 183454
rect 482902 183218 482904 183454
rect 482664 183134 482904 183218
rect 482664 182898 482666 183134
rect 482902 182898 482904 183134
rect 482664 182866 482904 182898
rect 491664 183454 491904 183486
rect 491664 183218 491666 183454
rect 491902 183218 491904 183454
rect 491664 183134 491904 183218
rect 491664 182898 491666 183134
rect 491902 182898 491904 183134
rect 491664 182866 491904 182898
rect 500664 183454 500904 183486
rect 500664 183218 500666 183454
rect 500902 183218 500904 183454
rect 500664 183134 500904 183218
rect 500664 182898 500666 183134
rect 500902 182898 500904 183134
rect 500664 182866 500904 182898
rect 509664 183454 509904 183486
rect 509664 183218 509666 183454
rect 509902 183218 509904 183454
rect 509664 183134 509904 183218
rect 509664 182898 509666 183134
rect 509902 182898 509904 183134
rect 509664 182866 509904 182898
rect 511466 183454 511706 183486
rect 511466 183218 511468 183454
rect 511704 183218 511706 183454
rect 511466 183134 511706 183218
rect 511466 182898 511468 183134
rect 511704 182898 511706 183134
rect 511466 182866 511706 182898
rect 512838 183454 513078 183486
rect 512838 183218 512840 183454
rect 513076 183218 513078 183454
rect 512838 183134 513078 183218
rect 512838 182898 512840 183134
rect 513076 182898 513078 183134
rect 512838 182866 513078 182898
rect 513684 183454 513924 183486
rect 513684 183218 513686 183454
rect 513922 183218 513924 183454
rect 513684 183134 513924 183218
rect 513684 182898 513686 183134
rect 513922 182898 513924 183134
rect 513684 182866 513924 182898
rect 522684 183454 522924 183486
rect 522684 183218 522686 183454
rect 522922 183218 522924 183454
rect 522684 183134 522924 183218
rect 522684 182898 522686 183134
rect 522922 182898 522924 183134
rect 522684 182866 522924 182898
rect 531684 183454 531924 183486
rect 531684 183218 531686 183454
rect 531922 183218 531924 183454
rect 531684 183134 531924 183218
rect 531684 182898 531686 183134
rect 531922 182898 531924 183134
rect 531684 182866 531924 182898
rect 540684 183454 540924 183486
rect 540684 183218 540686 183454
rect 540922 183218 540924 183454
rect 540684 183134 540924 183218
rect 540684 182898 540686 183134
rect 540922 182898 540924 183134
rect 540684 182866 540924 182898
rect 549684 183454 549924 183486
rect 549684 183218 549686 183454
rect 549922 183218 549924 183454
rect 549684 183134 549924 183218
rect 549684 182898 549686 183134
rect 549922 182898 549924 183134
rect 549684 182866 549924 182898
rect 551486 183454 551726 183486
rect 551486 183218 551488 183454
rect 551724 183218 551726 183454
rect 551486 183134 551726 183218
rect 551486 182898 551488 183134
rect 551724 182898 551726 183134
rect 551486 182866 551726 182898
rect 552858 183454 553098 183486
rect 552858 183218 552860 183454
rect 553096 183218 553098 183454
rect 552858 183134 553098 183218
rect 552858 182898 552860 183134
rect 553096 182898 553098 183134
rect 552858 182866 553098 182898
rect 553704 183454 553944 183486
rect 553704 183218 553706 183454
rect 553942 183218 553944 183454
rect 553704 183134 553944 183218
rect 553704 182898 553706 183134
rect 553942 182898 553944 183134
rect 553704 182866 553944 182898
rect 562704 183454 562944 183486
rect 562704 183218 562706 183454
rect 562942 183218 562944 183454
rect 562704 183134 562944 183218
rect 562704 182898 562706 183134
rect 562942 182898 562944 183134
rect 562704 182866 562944 182898
rect 571704 183454 571944 183486
rect 571704 183218 571706 183454
rect 571942 183218 571944 183454
rect 571704 183134 571944 183218
rect 571704 182898 571706 183134
rect 571942 182898 571944 183134
rect 571704 182866 571944 182898
rect 573474 183454 573714 183486
rect 573474 183218 573476 183454
rect 573712 183218 573714 183454
rect 573474 183134 573714 183218
rect 573474 182898 573476 183134
rect 573712 182898 573714 183134
rect 573474 182866 573714 182898
rect 578488 183454 579088 183486
rect 578488 183218 578670 183454
rect 578906 183218 579088 183454
rect 578488 183134 579088 183218
rect 578488 182898 578670 183134
rect 578906 182898 579088 183134
rect 578488 182866 579088 182898
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 4400 165454 5000 165486
rect 4400 165218 4582 165454
rect 4818 165218 5000 165454
rect 4400 165134 5000 165218
rect 4400 164898 4582 165134
rect 4818 164898 5000 165134
rect 4400 164866 5000 164898
rect 12230 165454 12470 165486
rect 12230 165218 12232 165454
rect 12468 165218 12470 165454
rect 12230 165134 12470 165218
rect 12230 164898 12232 165134
rect 12468 164898 12470 165134
rect 12230 164866 12470 164898
rect 13036 165454 13276 165486
rect 13036 165218 13038 165454
rect 13274 165218 13276 165454
rect 13036 165134 13276 165218
rect 13036 164898 13038 165134
rect 13274 164898 13276 165134
rect 13036 164866 13276 164898
rect 22036 165454 22276 165486
rect 22036 165218 22038 165454
rect 22274 165218 22276 165454
rect 22036 165134 22276 165218
rect 22036 164898 22038 165134
rect 22274 164898 22276 165134
rect 22036 164866 22276 164898
rect 27586 165454 27826 165486
rect 27586 165218 27588 165454
rect 27824 165218 27826 165454
rect 27586 165134 27826 165218
rect 27586 164898 27588 165134
rect 27824 164898 27826 165134
rect 27586 164866 27826 164898
rect 28238 165454 28478 165486
rect 28238 165218 28240 165454
rect 28476 165218 28478 165454
rect 28238 165134 28478 165218
rect 28238 164898 28240 165134
rect 28476 164898 28478 165134
rect 28238 164866 28478 164898
rect 29044 165454 29284 165486
rect 29044 165218 29046 165454
rect 29282 165218 29284 165454
rect 29044 165134 29284 165218
rect 29044 164898 29046 165134
rect 29282 164898 29284 165134
rect 29044 164866 29284 164898
rect 38044 165454 38284 165486
rect 38044 165218 38046 165454
rect 38282 165218 38284 165454
rect 38044 165134 38284 165218
rect 38044 164898 38046 165134
rect 38282 164898 38284 165134
rect 38044 164866 38284 164898
rect 47044 165454 47284 165486
rect 47044 165218 47046 165454
rect 47282 165218 47284 165454
rect 47044 165134 47284 165218
rect 47044 164898 47046 165134
rect 47282 164898 47284 165134
rect 47044 164866 47284 164898
rect 56044 165454 56284 165486
rect 56044 165218 56046 165454
rect 56282 165218 56284 165454
rect 56044 165134 56284 165218
rect 56044 164898 56046 165134
rect 56282 164898 56284 165134
rect 56044 164866 56284 164898
rect 65044 165454 65284 165486
rect 65044 165218 65046 165454
rect 65282 165218 65284 165454
rect 65044 165134 65284 165218
rect 65044 164898 65046 165134
rect 65282 164898 65284 165134
rect 65044 164866 65284 164898
rect 67606 165454 67846 165486
rect 67606 165218 67608 165454
rect 67844 165218 67846 165454
rect 67606 165134 67846 165218
rect 67606 164898 67608 165134
rect 67844 164898 67846 165134
rect 67606 164866 67846 164898
rect 68258 165454 68498 165486
rect 68258 165218 68260 165454
rect 68496 165218 68498 165454
rect 68258 165134 68498 165218
rect 68258 164898 68260 165134
rect 68496 164898 68498 165134
rect 68258 164866 68498 164898
rect 69064 165454 69304 165486
rect 69064 165218 69066 165454
rect 69302 165218 69304 165454
rect 69064 165134 69304 165218
rect 69064 164898 69066 165134
rect 69302 164898 69304 165134
rect 69064 164866 69304 164898
rect 78064 165454 78304 165486
rect 78064 165218 78066 165454
rect 78302 165218 78304 165454
rect 78064 165134 78304 165218
rect 78064 164898 78066 165134
rect 78302 164898 78304 165134
rect 78064 164866 78304 164898
rect 87064 165454 87304 165486
rect 87064 165218 87066 165454
rect 87302 165218 87304 165454
rect 87064 165134 87304 165218
rect 87064 164898 87066 165134
rect 87302 164898 87304 165134
rect 87064 164866 87304 164898
rect 96064 165454 96304 165486
rect 96064 165218 96066 165454
rect 96302 165218 96304 165454
rect 96064 165134 96304 165218
rect 96064 164898 96066 165134
rect 96302 164898 96304 165134
rect 96064 164866 96304 164898
rect 105064 165454 105304 165486
rect 105064 165218 105066 165454
rect 105302 165218 105304 165454
rect 105064 165134 105304 165218
rect 105064 164898 105066 165134
rect 105302 164898 105304 165134
rect 105064 164866 105304 164898
rect 107626 165454 107866 165486
rect 107626 165218 107628 165454
rect 107864 165218 107866 165454
rect 107626 165134 107866 165218
rect 107626 164898 107628 165134
rect 107864 164898 107866 165134
rect 107626 164866 107866 164898
rect 108278 165454 108518 165486
rect 108278 165218 108280 165454
rect 108516 165218 108518 165454
rect 108278 165134 108518 165218
rect 108278 164898 108280 165134
rect 108516 164898 108518 165134
rect 108278 164866 108518 164898
rect 109084 165454 109324 165486
rect 109084 165218 109086 165454
rect 109322 165218 109324 165454
rect 109084 165134 109324 165218
rect 109084 164898 109086 165134
rect 109322 164898 109324 165134
rect 109084 164866 109324 164898
rect 118084 165454 118324 165486
rect 118084 165218 118086 165454
rect 118322 165218 118324 165454
rect 118084 165134 118324 165218
rect 118084 164898 118086 165134
rect 118322 164898 118324 165134
rect 118084 164866 118324 164898
rect 127084 165454 127324 165486
rect 127084 165218 127086 165454
rect 127322 165218 127324 165454
rect 127084 165134 127324 165218
rect 127084 164898 127086 165134
rect 127322 164898 127324 165134
rect 127084 164866 127324 164898
rect 136084 165454 136324 165486
rect 136084 165218 136086 165454
rect 136322 165218 136324 165454
rect 136084 165134 136324 165218
rect 136084 164898 136086 165134
rect 136322 164898 136324 165134
rect 136084 164866 136324 164898
rect 145084 165454 145324 165486
rect 145084 165218 145086 165454
rect 145322 165218 145324 165454
rect 145084 165134 145324 165218
rect 145084 164898 145086 165134
rect 145322 164898 145324 165134
rect 145084 164866 145324 164898
rect 147646 165454 147886 165486
rect 147646 165218 147648 165454
rect 147884 165218 147886 165454
rect 147646 165134 147886 165218
rect 147646 164898 147648 165134
rect 147884 164898 147886 165134
rect 147646 164866 147886 164898
rect 149298 165454 149538 165486
rect 149298 165218 149300 165454
rect 149536 165218 149538 165454
rect 149298 165134 149538 165218
rect 149298 164898 149300 165134
rect 149536 164898 149538 165134
rect 149298 164866 149538 164898
rect 150104 165454 150344 165486
rect 150104 165218 150106 165454
rect 150342 165218 150344 165454
rect 150104 165134 150344 165218
rect 150104 164898 150106 165134
rect 150342 164898 150344 165134
rect 150104 164866 150344 164898
rect 159104 165454 159344 165486
rect 159104 165218 159106 165454
rect 159342 165218 159344 165454
rect 159104 165134 159344 165218
rect 159104 164898 159106 165134
rect 159342 164898 159344 165134
rect 159104 164866 159344 164898
rect 168104 165454 168344 165486
rect 168104 165218 168106 165454
rect 168342 165218 168344 165454
rect 168104 165134 168344 165218
rect 168104 164898 168106 165134
rect 168342 164898 168344 165134
rect 168104 164866 168344 164898
rect 177104 165454 177344 165486
rect 177104 165218 177106 165454
rect 177342 165218 177344 165454
rect 177104 165134 177344 165218
rect 177104 164898 177106 165134
rect 177342 164898 177344 165134
rect 177104 164866 177344 164898
rect 186104 165454 186344 165486
rect 186104 165218 186106 165454
rect 186342 165218 186344 165454
rect 186104 165134 186344 165218
rect 186104 164898 186106 165134
rect 186342 164898 186344 165134
rect 186104 164866 186344 164898
rect 188666 165454 188906 165486
rect 188666 165218 188668 165454
rect 188904 165218 188906 165454
rect 188666 165134 188906 165218
rect 188666 164898 188668 165134
rect 188904 164898 188906 165134
rect 188666 164866 188906 164898
rect 190318 165454 190558 165486
rect 190318 165218 190320 165454
rect 190556 165218 190558 165454
rect 190318 165134 190558 165218
rect 190318 164898 190320 165134
rect 190556 164898 190558 165134
rect 190318 164866 190558 164898
rect 191124 165454 191364 165486
rect 191124 165218 191126 165454
rect 191362 165218 191364 165454
rect 191124 165134 191364 165218
rect 191124 164898 191126 165134
rect 191362 164898 191364 165134
rect 191124 164866 191364 164898
rect 200124 165454 200364 165486
rect 200124 165218 200126 165454
rect 200362 165218 200364 165454
rect 200124 165134 200364 165218
rect 200124 164898 200126 165134
rect 200362 164898 200364 165134
rect 200124 164866 200364 164898
rect 209124 165454 209364 165486
rect 209124 165218 209126 165454
rect 209362 165218 209364 165454
rect 209124 165134 209364 165218
rect 209124 164898 209126 165134
rect 209362 164898 209364 165134
rect 209124 164866 209364 164898
rect 218124 165454 218364 165486
rect 218124 165218 218126 165454
rect 218362 165218 218364 165454
rect 218124 165134 218364 165218
rect 218124 164898 218126 165134
rect 218362 164898 218364 165134
rect 218124 164866 218364 164898
rect 227124 165454 227364 165486
rect 227124 165218 227126 165454
rect 227362 165218 227364 165454
rect 227124 165134 227364 165218
rect 227124 164898 227126 165134
rect 227362 164898 227364 165134
rect 227124 164866 227364 164898
rect 229686 165454 229926 165486
rect 229686 165218 229688 165454
rect 229924 165218 229926 165454
rect 229686 165134 229926 165218
rect 229686 164898 229688 165134
rect 229924 164898 229926 165134
rect 229686 164866 229926 164898
rect 230338 165454 230578 165486
rect 230338 165218 230340 165454
rect 230576 165218 230578 165454
rect 230338 165134 230578 165218
rect 230338 164898 230340 165134
rect 230576 164898 230578 165134
rect 230338 164866 230578 164898
rect 231144 165454 231384 165486
rect 231144 165218 231146 165454
rect 231382 165218 231384 165454
rect 231144 165134 231384 165218
rect 231144 164898 231146 165134
rect 231382 164898 231384 165134
rect 231144 164866 231384 164898
rect 240144 165454 240384 165486
rect 240144 165218 240146 165454
rect 240382 165218 240384 165454
rect 240144 165134 240384 165218
rect 240144 164898 240146 165134
rect 240382 164898 240384 165134
rect 240144 164866 240384 164898
rect 249144 165454 249384 165486
rect 249144 165218 249146 165454
rect 249382 165218 249384 165454
rect 249144 165134 249384 165218
rect 249144 164898 249146 165134
rect 249382 164898 249384 165134
rect 249144 164866 249384 164898
rect 258144 165454 258384 165486
rect 258144 165218 258146 165454
rect 258382 165218 258384 165454
rect 258144 165134 258384 165218
rect 258144 164898 258146 165134
rect 258382 164898 258384 165134
rect 258144 164866 258384 164898
rect 267144 165454 267384 165486
rect 267144 165218 267146 165454
rect 267382 165218 267384 165454
rect 267144 165134 267384 165218
rect 267144 164898 267146 165134
rect 267382 164898 267384 165134
rect 267144 164866 267384 164898
rect 269706 165454 269946 165486
rect 269706 165218 269708 165454
rect 269944 165218 269946 165454
rect 269706 165134 269946 165218
rect 269706 164898 269708 165134
rect 269944 164898 269946 165134
rect 269706 164866 269946 164898
rect 270358 165454 270598 165486
rect 270358 165218 270360 165454
rect 270596 165218 270598 165454
rect 270358 165134 270598 165218
rect 270358 164898 270360 165134
rect 270596 164898 270598 165134
rect 270358 164866 270598 164898
rect 271164 165454 271404 165486
rect 271164 165218 271166 165454
rect 271402 165218 271404 165454
rect 271164 165134 271404 165218
rect 271164 164898 271166 165134
rect 271402 164898 271404 165134
rect 271164 164866 271404 164898
rect 280164 165454 280404 165486
rect 280164 165218 280166 165454
rect 280402 165218 280404 165454
rect 280164 165134 280404 165218
rect 280164 164898 280166 165134
rect 280402 164898 280404 165134
rect 280164 164866 280404 164898
rect 289164 165454 289404 165486
rect 289164 165218 289166 165454
rect 289402 165218 289404 165454
rect 289164 165134 289404 165218
rect 289164 164898 289166 165134
rect 289402 164898 289404 165134
rect 289164 164866 289404 164898
rect 298164 165454 298404 165486
rect 298164 165218 298166 165454
rect 298402 165218 298404 165454
rect 298164 165134 298404 165218
rect 298164 164898 298166 165134
rect 298402 164898 298404 165134
rect 298164 164866 298404 164898
rect 307164 165454 307404 165486
rect 307164 165218 307166 165454
rect 307402 165218 307404 165454
rect 307164 165134 307404 165218
rect 307164 164898 307166 165134
rect 307402 164898 307404 165134
rect 307164 164866 307404 164898
rect 309726 165454 309966 165486
rect 309726 165218 309728 165454
rect 309964 165218 309966 165454
rect 309726 165134 309966 165218
rect 309726 164898 309728 165134
rect 309964 164898 309966 165134
rect 309726 164866 309966 164898
rect 311378 165454 311618 165486
rect 311378 165218 311380 165454
rect 311616 165218 311618 165454
rect 311378 165134 311618 165218
rect 311378 164898 311380 165134
rect 311616 164898 311618 165134
rect 311378 164866 311618 164898
rect 312184 165454 312424 165486
rect 312184 165218 312186 165454
rect 312422 165218 312424 165454
rect 312184 165134 312424 165218
rect 312184 164898 312186 165134
rect 312422 164898 312424 165134
rect 312184 164866 312424 164898
rect 321184 165454 321424 165486
rect 321184 165218 321186 165454
rect 321422 165218 321424 165454
rect 321184 165134 321424 165218
rect 321184 164898 321186 165134
rect 321422 164898 321424 165134
rect 321184 164866 321424 164898
rect 330184 165454 330424 165486
rect 330184 165218 330186 165454
rect 330422 165218 330424 165454
rect 330184 165134 330424 165218
rect 330184 164898 330186 165134
rect 330422 164898 330424 165134
rect 330184 164866 330424 164898
rect 339184 165454 339424 165486
rect 339184 165218 339186 165454
rect 339422 165218 339424 165454
rect 339184 165134 339424 165218
rect 339184 164898 339186 165134
rect 339422 164898 339424 165134
rect 339184 164866 339424 164898
rect 348184 165454 348424 165486
rect 348184 165218 348186 165454
rect 348422 165218 348424 165454
rect 348184 165134 348424 165218
rect 348184 164898 348186 165134
rect 348422 164898 348424 165134
rect 348184 164866 348424 164898
rect 350746 165454 350986 165486
rect 350746 165218 350748 165454
rect 350984 165218 350986 165454
rect 350746 165134 350986 165218
rect 350746 164898 350748 165134
rect 350984 164898 350986 165134
rect 350746 164866 350986 164898
rect 352398 165454 352638 165486
rect 352398 165218 352400 165454
rect 352636 165218 352638 165454
rect 352398 165134 352638 165218
rect 352398 164898 352400 165134
rect 352636 164898 352638 165134
rect 352398 164866 352638 164898
rect 353204 165454 353444 165486
rect 353204 165218 353206 165454
rect 353442 165218 353444 165454
rect 353204 165134 353444 165218
rect 353204 164898 353206 165134
rect 353442 164898 353444 165134
rect 353204 164866 353444 164898
rect 362204 165454 362444 165486
rect 362204 165218 362206 165454
rect 362442 165218 362444 165454
rect 362204 165134 362444 165218
rect 362204 164898 362206 165134
rect 362442 164898 362444 165134
rect 362204 164866 362444 164898
rect 371204 165454 371444 165486
rect 371204 165218 371206 165454
rect 371442 165218 371444 165454
rect 371204 165134 371444 165218
rect 371204 164898 371206 165134
rect 371442 164898 371444 165134
rect 371204 164866 371444 164898
rect 380204 165454 380444 165486
rect 380204 165218 380206 165454
rect 380442 165218 380444 165454
rect 380204 165134 380444 165218
rect 380204 164898 380206 165134
rect 380442 164898 380444 165134
rect 380204 164866 380444 164898
rect 389204 165454 389444 165486
rect 389204 165218 389206 165454
rect 389442 165218 389444 165454
rect 389204 165134 389444 165218
rect 389204 164898 389206 165134
rect 389442 164898 389444 165134
rect 389204 164866 389444 164898
rect 391766 165454 392006 165486
rect 391766 165218 391768 165454
rect 392004 165218 392006 165454
rect 391766 165134 392006 165218
rect 391766 164898 391768 165134
rect 392004 164898 392006 165134
rect 391766 164866 392006 164898
rect 392418 165454 392658 165486
rect 392418 165218 392420 165454
rect 392656 165218 392658 165454
rect 392418 165134 392658 165218
rect 392418 164898 392420 165134
rect 392656 164898 392658 165134
rect 392418 164866 392658 164898
rect 393224 165454 393464 165486
rect 393224 165218 393226 165454
rect 393462 165218 393464 165454
rect 393224 165134 393464 165218
rect 393224 164898 393226 165134
rect 393462 164898 393464 165134
rect 393224 164866 393464 164898
rect 402224 165454 402464 165486
rect 402224 165218 402226 165454
rect 402462 165218 402464 165454
rect 402224 165134 402464 165218
rect 402224 164898 402226 165134
rect 402462 164898 402464 165134
rect 402224 164866 402464 164898
rect 411224 165454 411464 165486
rect 411224 165218 411226 165454
rect 411462 165218 411464 165454
rect 411224 165134 411464 165218
rect 411224 164898 411226 165134
rect 411462 164898 411464 165134
rect 411224 164866 411464 164898
rect 420224 165454 420464 165486
rect 420224 165218 420226 165454
rect 420462 165218 420464 165454
rect 420224 165134 420464 165218
rect 420224 164898 420226 165134
rect 420462 164898 420464 165134
rect 420224 164866 420464 164898
rect 429224 165454 429464 165486
rect 429224 165218 429226 165454
rect 429462 165218 429464 165454
rect 429224 165134 429464 165218
rect 429224 164898 429226 165134
rect 429462 164898 429464 165134
rect 429224 164866 429464 164898
rect 431786 165454 432026 165486
rect 431786 165218 431788 165454
rect 432024 165218 432026 165454
rect 431786 165134 432026 165218
rect 431786 164898 431788 165134
rect 432024 164898 432026 165134
rect 431786 164866 432026 164898
rect 432438 165454 432678 165486
rect 432438 165218 432440 165454
rect 432676 165218 432678 165454
rect 432438 165134 432678 165218
rect 432438 164898 432440 165134
rect 432676 164898 432678 165134
rect 432438 164866 432678 164898
rect 433244 165454 433484 165486
rect 433244 165218 433246 165454
rect 433482 165218 433484 165454
rect 433244 165134 433484 165218
rect 433244 164898 433246 165134
rect 433482 164898 433484 165134
rect 433244 164866 433484 164898
rect 442244 165454 442484 165486
rect 442244 165218 442246 165454
rect 442482 165218 442484 165454
rect 442244 165134 442484 165218
rect 442244 164898 442246 165134
rect 442482 164898 442484 165134
rect 442244 164866 442484 164898
rect 451244 165454 451484 165486
rect 451244 165218 451246 165454
rect 451482 165218 451484 165454
rect 451244 165134 451484 165218
rect 451244 164898 451246 165134
rect 451482 164898 451484 165134
rect 451244 164866 451484 164898
rect 460244 165454 460484 165486
rect 460244 165218 460246 165454
rect 460482 165218 460484 165454
rect 460244 165134 460484 165218
rect 460244 164898 460246 165134
rect 460482 164898 460484 165134
rect 460244 164866 460484 164898
rect 469244 165454 469484 165486
rect 469244 165218 469246 165454
rect 469482 165218 469484 165454
rect 469244 165134 469484 165218
rect 469244 164898 469246 165134
rect 469482 164898 469484 165134
rect 469244 164866 469484 164898
rect 471806 165454 472046 165486
rect 471806 165218 471808 165454
rect 472044 165218 472046 165454
rect 471806 165134 472046 165218
rect 471806 164898 471808 165134
rect 472044 164898 472046 165134
rect 471806 164866 472046 164898
rect 472458 165454 472698 165486
rect 472458 165218 472460 165454
rect 472696 165218 472698 165454
rect 472458 165134 472698 165218
rect 472458 164898 472460 165134
rect 472696 164898 472698 165134
rect 472458 164866 472698 164898
rect 473264 165454 473504 165486
rect 473264 165218 473266 165454
rect 473502 165218 473504 165454
rect 473264 165134 473504 165218
rect 473264 164898 473266 165134
rect 473502 164898 473504 165134
rect 473264 164866 473504 164898
rect 482264 165454 482504 165486
rect 482264 165218 482266 165454
rect 482502 165218 482504 165454
rect 482264 165134 482504 165218
rect 482264 164898 482266 165134
rect 482502 164898 482504 165134
rect 482264 164866 482504 164898
rect 491264 165454 491504 165486
rect 491264 165218 491266 165454
rect 491502 165218 491504 165454
rect 491264 165134 491504 165218
rect 491264 164898 491266 165134
rect 491502 164898 491504 165134
rect 491264 164866 491504 164898
rect 500264 165454 500504 165486
rect 500264 165218 500266 165454
rect 500502 165218 500504 165454
rect 500264 165134 500504 165218
rect 500264 164898 500266 165134
rect 500502 164898 500504 165134
rect 500264 164866 500504 164898
rect 509264 165454 509504 165486
rect 509264 165218 509266 165454
rect 509502 165218 509504 165454
rect 509264 165134 509504 165218
rect 509264 164898 509266 165134
rect 509502 164898 509504 165134
rect 509264 164866 509504 164898
rect 511826 165454 512066 165486
rect 511826 165218 511828 165454
rect 512064 165218 512066 165454
rect 511826 165134 512066 165218
rect 511826 164898 511828 165134
rect 512064 164898 512066 165134
rect 511826 164866 512066 164898
rect 512478 165454 512718 165486
rect 512478 165218 512480 165454
rect 512716 165218 512718 165454
rect 512478 165134 512718 165218
rect 512478 164898 512480 165134
rect 512716 164898 512718 165134
rect 512478 164866 512718 164898
rect 513284 165454 513524 165486
rect 513284 165218 513286 165454
rect 513522 165218 513524 165454
rect 513284 165134 513524 165218
rect 513284 164898 513286 165134
rect 513522 164898 513524 165134
rect 513284 164866 513524 164898
rect 522284 165454 522524 165486
rect 522284 165218 522286 165454
rect 522522 165218 522524 165454
rect 522284 165134 522524 165218
rect 522284 164898 522286 165134
rect 522522 164898 522524 165134
rect 522284 164866 522524 164898
rect 531284 165454 531524 165486
rect 531284 165218 531286 165454
rect 531522 165218 531524 165454
rect 531284 165134 531524 165218
rect 531284 164898 531286 165134
rect 531522 164898 531524 165134
rect 531284 164866 531524 164898
rect 540284 165454 540524 165486
rect 540284 165218 540286 165454
rect 540522 165218 540524 165454
rect 540284 165134 540524 165218
rect 540284 164898 540286 165134
rect 540522 164898 540524 165134
rect 540284 164866 540524 164898
rect 549284 165454 549524 165486
rect 549284 165218 549286 165454
rect 549522 165218 549524 165454
rect 549284 165134 549524 165218
rect 549284 164898 549286 165134
rect 549522 164898 549524 165134
rect 549284 164866 549524 164898
rect 551846 165454 552086 165486
rect 551846 165218 551848 165454
rect 552084 165218 552086 165454
rect 551846 165134 552086 165218
rect 551846 164898 551848 165134
rect 552084 164898 552086 165134
rect 551846 164866 552086 164898
rect 552498 165454 552738 165486
rect 552498 165218 552500 165454
rect 552736 165218 552738 165454
rect 552498 165134 552738 165218
rect 552498 164898 552500 165134
rect 552736 164898 552738 165134
rect 552498 164866 552738 164898
rect 553304 165454 553544 165486
rect 553304 165218 553306 165454
rect 553542 165218 553544 165454
rect 553304 165134 553544 165218
rect 553304 164898 553306 165134
rect 553542 164898 553544 165134
rect 553304 164866 553544 164898
rect 562304 165454 562544 165486
rect 562304 165218 562306 165454
rect 562542 165218 562544 165454
rect 562304 165134 562544 165218
rect 562304 164898 562306 165134
rect 562542 164898 562544 165134
rect 562304 164866 562544 164898
rect 571304 165454 571544 165486
rect 571304 165218 571306 165454
rect 571542 165218 571544 165454
rect 571304 165134 571544 165218
rect 571304 164898 571306 165134
rect 571542 164898 571544 165134
rect 571304 164866 571544 164898
rect 573834 165454 574074 165486
rect 573834 165218 573836 165454
rect 574072 165218 574074 165454
rect 573834 165134 574074 165218
rect 573834 164898 573836 165134
rect 574072 164898 574074 165134
rect 573834 164866 574074 164898
rect 579288 165454 579888 165486
rect 579288 165218 579470 165454
rect 579706 165218 579888 165454
rect 579288 165134 579888 165218
rect 579288 164898 579470 165134
rect 579706 164898 579888 165134
rect 579288 164866 579888 164898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect 5200 147454 5800 147486
rect 5200 147218 5382 147454
rect 5618 147218 5800 147454
rect 5200 147134 5800 147218
rect 5200 146898 5382 147134
rect 5618 146898 5800 147134
rect 5200 146866 5800 146898
rect 12590 147454 12830 147486
rect 12590 147218 12592 147454
rect 12828 147218 12830 147454
rect 12590 147134 12830 147218
rect 12590 146898 12592 147134
rect 12828 146898 12830 147134
rect 12590 146866 12830 146898
rect 13436 147454 13676 147486
rect 13436 147218 13438 147454
rect 13674 147218 13676 147454
rect 13436 147134 13676 147218
rect 13436 146898 13438 147134
rect 13674 146898 13676 147134
rect 13436 146866 13676 146898
rect 22436 147454 22676 147486
rect 22436 147218 22438 147454
rect 22674 147218 22676 147454
rect 22436 147134 22676 147218
rect 22436 146898 22438 147134
rect 22674 146898 22676 147134
rect 22436 146866 22676 146898
rect 27226 147454 27466 147486
rect 27226 147218 27228 147454
rect 27464 147218 27466 147454
rect 27226 147134 27466 147218
rect 27226 146898 27228 147134
rect 27464 146898 27466 147134
rect 27226 146866 27466 146898
rect 28598 147454 28838 147486
rect 28598 147218 28600 147454
rect 28836 147218 28838 147454
rect 28598 147134 28838 147218
rect 28598 146898 28600 147134
rect 28836 146898 28838 147134
rect 28598 146866 28838 146898
rect 29444 147454 29684 147486
rect 29444 147218 29446 147454
rect 29682 147218 29684 147454
rect 29444 147134 29684 147218
rect 29444 146898 29446 147134
rect 29682 146898 29684 147134
rect 29444 146866 29684 146898
rect 38444 147454 38684 147486
rect 38444 147218 38446 147454
rect 38682 147218 38684 147454
rect 38444 147134 38684 147218
rect 38444 146898 38446 147134
rect 38682 146898 38684 147134
rect 38444 146866 38684 146898
rect 47444 147454 47684 147486
rect 47444 147218 47446 147454
rect 47682 147218 47684 147454
rect 47444 147134 47684 147218
rect 47444 146898 47446 147134
rect 47682 146898 47684 147134
rect 47444 146866 47684 146898
rect 56444 147454 56684 147486
rect 56444 147218 56446 147454
rect 56682 147218 56684 147454
rect 56444 147134 56684 147218
rect 56444 146898 56446 147134
rect 56682 146898 56684 147134
rect 56444 146866 56684 146898
rect 65444 147454 65684 147486
rect 65444 147218 65446 147454
rect 65682 147218 65684 147454
rect 65444 147134 65684 147218
rect 65444 146898 65446 147134
rect 65682 146898 65684 147134
rect 65444 146866 65684 146898
rect 67246 147454 67486 147486
rect 67246 147218 67248 147454
rect 67484 147218 67486 147454
rect 67246 147134 67486 147218
rect 67246 146898 67248 147134
rect 67484 146898 67486 147134
rect 67246 146866 67486 146898
rect 68618 147454 68858 147486
rect 68618 147218 68620 147454
rect 68856 147218 68858 147454
rect 68618 147134 68858 147218
rect 68618 146898 68620 147134
rect 68856 146898 68858 147134
rect 68618 146866 68858 146898
rect 69464 147454 69704 147486
rect 69464 147218 69466 147454
rect 69702 147218 69704 147454
rect 69464 147134 69704 147218
rect 69464 146898 69466 147134
rect 69702 146898 69704 147134
rect 69464 146866 69704 146898
rect 78464 147454 78704 147486
rect 78464 147218 78466 147454
rect 78702 147218 78704 147454
rect 78464 147134 78704 147218
rect 78464 146898 78466 147134
rect 78702 146898 78704 147134
rect 78464 146866 78704 146898
rect 87464 147454 87704 147486
rect 87464 147218 87466 147454
rect 87702 147218 87704 147454
rect 87464 147134 87704 147218
rect 87464 146898 87466 147134
rect 87702 146898 87704 147134
rect 87464 146866 87704 146898
rect 96464 147454 96704 147486
rect 96464 147218 96466 147454
rect 96702 147218 96704 147454
rect 96464 147134 96704 147218
rect 96464 146898 96466 147134
rect 96702 146898 96704 147134
rect 96464 146866 96704 146898
rect 105464 147454 105704 147486
rect 105464 147218 105466 147454
rect 105702 147218 105704 147454
rect 105464 147134 105704 147218
rect 105464 146898 105466 147134
rect 105702 146898 105704 147134
rect 105464 146866 105704 146898
rect 107266 147454 107506 147486
rect 107266 147218 107268 147454
rect 107504 147218 107506 147454
rect 107266 147134 107506 147218
rect 107266 146898 107268 147134
rect 107504 146898 107506 147134
rect 107266 146866 107506 146898
rect 108638 147454 108878 147486
rect 108638 147218 108640 147454
rect 108876 147218 108878 147454
rect 108638 147134 108878 147218
rect 108638 146898 108640 147134
rect 108876 146898 108878 147134
rect 108638 146866 108878 146898
rect 109484 147454 109724 147486
rect 109484 147218 109486 147454
rect 109722 147218 109724 147454
rect 109484 147134 109724 147218
rect 109484 146898 109486 147134
rect 109722 146898 109724 147134
rect 109484 146866 109724 146898
rect 118484 147454 118724 147486
rect 118484 147218 118486 147454
rect 118722 147218 118724 147454
rect 118484 147134 118724 147218
rect 118484 146898 118486 147134
rect 118722 146898 118724 147134
rect 118484 146866 118724 146898
rect 127484 147454 127724 147486
rect 127484 147218 127486 147454
rect 127722 147218 127724 147454
rect 127484 147134 127724 147218
rect 127484 146898 127486 147134
rect 127722 146898 127724 147134
rect 127484 146866 127724 146898
rect 136484 147454 136724 147486
rect 136484 147218 136486 147454
rect 136722 147218 136724 147454
rect 136484 147134 136724 147218
rect 136484 146898 136486 147134
rect 136722 146898 136724 147134
rect 136484 146866 136724 146898
rect 145484 147454 145724 147486
rect 145484 147218 145486 147454
rect 145722 147218 145724 147454
rect 145484 147134 145724 147218
rect 145484 146898 145486 147134
rect 145722 146898 145724 147134
rect 145484 146866 145724 146898
rect 147286 147454 147526 147486
rect 147286 147218 147288 147454
rect 147524 147218 147526 147454
rect 147286 147134 147526 147218
rect 147286 146898 147288 147134
rect 147524 146898 147526 147134
rect 147286 146866 147526 146898
rect 149658 147454 149898 147486
rect 149658 147218 149660 147454
rect 149896 147218 149898 147454
rect 149658 147134 149898 147218
rect 149658 146898 149660 147134
rect 149896 146898 149898 147134
rect 149658 146866 149898 146898
rect 150504 147454 150744 147486
rect 150504 147218 150506 147454
rect 150742 147218 150744 147454
rect 150504 147134 150744 147218
rect 150504 146898 150506 147134
rect 150742 146898 150744 147134
rect 150504 146866 150744 146898
rect 159504 147454 159744 147486
rect 159504 147218 159506 147454
rect 159742 147218 159744 147454
rect 159504 147134 159744 147218
rect 159504 146898 159506 147134
rect 159742 146898 159744 147134
rect 159504 146866 159744 146898
rect 168504 147454 168744 147486
rect 168504 147218 168506 147454
rect 168742 147218 168744 147454
rect 168504 147134 168744 147218
rect 168504 146898 168506 147134
rect 168742 146898 168744 147134
rect 168504 146866 168744 146898
rect 177504 147454 177744 147486
rect 177504 147218 177506 147454
rect 177742 147218 177744 147454
rect 177504 147134 177744 147218
rect 177504 146898 177506 147134
rect 177742 146898 177744 147134
rect 177504 146866 177744 146898
rect 186504 147454 186744 147486
rect 186504 147218 186506 147454
rect 186742 147218 186744 147454
rect 186504 147134 186744 147218
rect 186504 146898 186506 147134
rect 186742 146898 186744 147134
rect 186504 146866 186744 146898
rect 188306 147454 188546 147486
rect 188306 147218 188308 147454
rect 188544 147218 188546 147454
rect 188306 147134 188546 147218
rect 188306 146898 188308 147134
rect 188544 146898 188546 147134
rect 188306 146866 188546 146898
rect 190678 147454 190918 147486
rect 190678 147218 190680 147454
rect 190916 147218 190918 147454
rect 190678 147134 190918 147218
rect 190678 146898 190680 147134
rect 190916 146898 190918 147134
rect 190678 146866 190918 146898
rect 191524 147454 191764 147486
rect 191524 147218 191526 147454
rect 191762 147218 191764 147454
rect 191524 147134 191764 147218
rect 191524 146898 191526 147134
rect 191762 146898 191764 147134
rect 191524 146866 191764 146898
rect 200524 147454 200764 147486
rect 200524 147218 200526 147454
rect 200762 147218 200764 147454
rect 200524 147134 200764 147218
rect 200524 146898 200526 147134
rect 200762 146898 200764 147134
rect 200524 146866 200764 146898
rect 209524 147454 209764 147486
rect 209524 147218 209526 147454
rect 209762 147218 209764 147454
rect 209524 147134 209764 147218
rect 209524 146898 209526 147134
rect 209762 146898 209764 147134
rect 209524 146866 209764 146898
rect 218524 147454 218764 147486
rect 218524 147218 218526 147454
rect 218762 147218 218764 147454
rect 218524 147134 218764 147218
rect 218524 146898 218526 147134
rect 218762 146898 218764 147134
rect 218524 146866 218764 146898
rect 227524 147454 227764 147486
rect 227524 147218 227526 147454
rect 227762 147218 227764 147454
rect 227524 147134 227764 147218
rect 227524 146898 227526 147134
rect 227762 146898 227764 147134
rect 227524 146866 227764 146898
rect 229326 147454 229566 147486
rect 229326 147218 229328 147454
rect 229564 147218 229566 147454
rect 229326 147134 229566 147218
rect 229326 146898 229328 147134
rect 229564 146898 229566 147134
rect 229326 146866 229566 146898
rect 230698 147454 230938 147486
rect 230698 147218 230700 147454
rect 230936 147218 230938 147454
rect 230698 147134 230938 147218
rect 230698 146898 230700 147134
rect 230936 146898 230938 147134
rect 230698 146866 230938 146898
rect 231544 147454 231784 147486
rect 231544 147218 231546 147454
rect 231782 147218 231784 147454
rect 231544 147134 231784 147218
rect 231544 146898 231546 147134
rect 231782 146898 231784 147134
rect 231544 146866 231784 146898
rect 240544 147454 240784 147486
rect 240544 147218 240546 147454
rect 240782 147218 240784 147454
rect 240544 147134 240784 147218
rect 240544 146898 240546 147134
rect 240782 146898 240784 147134
rect 240544 146866 240784 146898
rect 249544 147454 249784 147486
rect 249544 147218 249546 147454
rect 249782 147218 249784 147454
rect 249544 147134 249784 147218
rect 249544 146898 249546 147134
rect 249782 146898 249784 147134
rect 249544 146866 249784 146898
rect 258544 147454 258784 147486
rect 258544 147218 258546 147454
rect 258782 147218 258784 147454
rect 258544 147134 258784 147218
rect 258544 146898 258546 147134
rect 258782 146898 258784 147134
rect 258544 146866 258784 146898
rect 267544 147454 267784 147486
rect 267544 147218 267546 147454
rect 267782 147218 267784 147454
rect 267544 147134 267784 147218
rect 267544 146898 267546 147134
rect 267782 146898 267784 147134
rect 267544 146866 267784 146898
rect 269346 147454 269586 147486
rect 269346 147218 269348 147454
rect 269584 147218 269586 147454
rect 269346 147134 269586 147218
rect 269346 146898 269348 147134
rect 269584 146898 269586 147134
rect 269346 146866 269586 146898
rect 270718 147454 270958 147486
rect 270718 147218 270720 147454
rect 270956 147218 270958 147454
rect 270718 147134 270958 147218
rect 270718 146898 270720 147134
rect 270956 146898 270958 147134
rect 270718 146866 270958 146898
rect 271564 147454 271804 147486
rect 271564 147218 271566 147454
rect 271802 147218 271804 147454
rect 271564 147134 271804 147218
rect 271564 146898 271566 147134
rect 271802 146898 271804 147134
rect 271564 146866 271804 146898
rect 280564 147454 280804 147486
rect 280564 147218 280566 147454
rect 280802 147218 280804 147454
rect 280564 147134 280804 147218
rect 280564 146898 280566 147134
rect 280802 146898 280804 147134
rect 280564 146866 280804 146898
rect 289564 147454 289804 147486
rect 289564 147218 289566 147454
rect 289802 147218 289804 147454
rect 289564 147134 289804 147218
rect 289564 146898 289566 147134
rect 289802 146898 289804 147134
rect 289564 146866 289804 146898
rect 298564 147454 298804 147486
rect 298564 147218 298566 147454
rect 298802 147218 298804 147454
rect 298564 147134 298804 147218
rect 298564 146898 298566 147134
rect 298802 146898 298804 147134
rect 298564 146866 298804 146898
rect 307564 147454 307804 147486
rect 307564 147218 307566 147454
rect 307802 147218 307804 147454
rect 307564 147134 307804 147218
rect 307564 146898 307566 147134
rect 307802 146898 307804 147134
rect 307564 146866 307804 146898
rect 309366 147454 309606 147486
rect 309366 147218 309368 147454
rect 309604 147218 309606 147454
rect 309366 147134 309606 147218
rect 309366 146898 309368 147134
rect 309604 146898 309606 147134
rect 309366 146866 309606 146898
rect 311738 147454 311978 147486
rect 311738 147218 311740 147454
rect 311976 147218 311978 147454
rect 311738 147134 311978 147218
rect 311738 146898 311740 147134
rect 311976 146898 311978 147134
rect 311738 146866 311978 146898
rect 312584 147454 312824 147486
rect 312584 147218 312586 147454
rect 312822 147218 312824 147454
rect 312584 147134 312824 147218
rect 312584 146898 312586 147134
rect 312822 146898 312824 147134
rect 312584 146866 312824 146898
rect 321584 147454 321824 147486
rect 321584 147218 321586 147454
rect 321822 147218 321824 147454
rect 321584 147134 321824 147218
rect 321584 146898 321586 147134
rect 321822 146898 321824 147134
rect 321584 146866 321824 146898
rect 330584 147454 330824 147486
rect 330584 147218 330586 147454
rect 330822 147218 330824 147454
rect 330584 147134 330824 147218
rect 330584 146898 330586 147134
rect 330822 146898 330824 147134
rect 330584 146866 330824 146898
rect 339584 147454 339824 147486
rect 339584 147218 339586 147454
rect 339822 147218 339824 147454
rect 339584 147134 339824 147218
rect 339584 146898 339586 147134
rect 339822 146898 339824 147134
rect 339584 146866 339824 146898
rect 348584 147454 348824 147486
rect 348584 147218 348586 147454
rect 348822 147218 348824 147454
rect 348584 147134 348824 147218
rect 348584 146898 348586 147134
rect 348822 146898 348824 147134
rect 348584 146866 348824 146898
rect 350386 147454 350626 147486
rect 350386 147218 350388 147454
rect 350624 147218 350626 147454
rect 350386 147134 350626 147218
rect 350386 146898 350388 147134
rect 350624 146898 350626 147134
rect 350386 146866 350626 146898
rect 352758 147454 352998 147486
rect 352758 147218 352760 147454
rect 352996 147218 352998 147454
rect 352758 147134 352998 147218
rect 352758 146898 352760 147134
rect 352996 146898 352998 147134
rect 352758 146866 352998 146898
rect 353604 147454 353844 147486
rect 353604 147218 353606 147454
rect 353842 147218 353844 147454
rect 353604 147134 353844 147218
rect 353604 146898 353606 147134
rect 353842 146898 353844 147134
rect 353604 146866 353844 146898
rect 362604 147454 362844 147486
rect 362604 147218 362606 147454
rect 362842 147218 362844 147454
rect 362604 147134 362844 147218
rect 362604 146898 362606 147134
rect 362842 146898 362844 147134
rect 362604 146866 362844 146898
rect 371604 147454 371844 147486
rect 371604 147218 371606 147454
rect 371842 147218 371844 147454
rect 371604 147134 371844 147218
rect 371604 146898 371606 147134
rect 371842 146898 371844 147134
rect 371604 146866 371844 146898
rect 380604 147454 380844 147486
rect 380604 147218 380606 147454
rect 380842 147218 380844 147454
rect 380604 147134 380844 147218
rect 380604 146898 380606 147134
rect 380842 146898 380844 147134
rect 380604 146866 380844 146898
rect 389604 147454 389844 147486
rect 389604 147218 389606 147454
rect 389842 147218 389844 147454
rect 389604 147134 389844 147218
rect 389604 146898 389606 147134
rect 389842 146898 389844 147134
rect 389604 146866 389844 146898
rect 391406 147454 391646 147486
rect 391406 147218 391408 147454
rect 391644 147218 391646 147454
rect 391406 147134 391646 147218
rect 391406 146898 391408 147134
rect 391644 146898 391646 147134
rect 391406 146866 391646 146898
rect 392778 147454 393018 147486
rect 392778 147218 392780 147454
rect 393016 147218 393018 147454
rect 392778 147134 393018 147218
rect 392778 146898 392780 147134
rect 393016 146898 393018 147134
rect 392778 146866 393018 146898
rect 393624 147454 393864 147486
rect 393624 147218 393626 147454
rect 393862 147218 393864 147454
rect 393624 147134 393864 147218
rect 393624 146898 393626 147134
rect 393862 146898 393864 147134
rect 393624 146866 393864 146898
rect 402624 147454 402864 147486
rect 402624 147218 402626 147454
rect 402862 147218 402864 147454
rect 402624 147134 402864 147218
rect 402624 146898 402626 147134
rect 402862 146898 402864 147134
rect 402624 146866 402864 146898
rect 411624 147454 411864 147486
rect 411624 147218 411626 147454
rect 411862 147218 411864 147454
rect 411624 147134 411864 147218
rect 411624 146898 411626 147134
rect 411862 146898 411864 147134
rect 411624 146866 411864 146898
rect 420624 147454 420864 147486
rect 420624 147218 420626 147454
rect 420862 147218 420864 147454
rect 420624 147134 420864 147218
rect 420624 146898 420626 147134
rect 420862 146898 420864 147134
rect 420624 146866 420864 146898
rect 429624 147454 429864 147486
rect 429624 147218 429626 147454
rect 429862 147218 429864 147454
rect 429624 147134 429864 147218
rect 429624 146898 429626 147134
rect 429862 146898 429864 147134
rect 429624 146866 429864 146898
rect 431426 147454 431666 147486
rect 431426 147218 431428 147454
rect 431664 147218 431666 147454
rect 431426 147134 431666 147218
rect 431426 146898 431428 147134
rect 431664 146898 431666 147134
rect 431426 146866 431666 146898
rect 432798 147454 433038 147486
rect 432798 147218 432800 147454
rect 433036 147218 433038 147454
rect 432798 147134 433038 147218
rect 432798 146898 432800 147134
rect 433036 146898 433038 147134
rect 432798 146866 433038 146898
rect 433644 147454 433884 147486
rect 433644 147218 433646 147454
rect 433882 147218 433884 147454
rect 433644 147134 433884 147218
rect 433644 146898 433646 147134
rect 433882 146898 433884 147134
rect 433644 146866 433884 146898
rect 442644 147454 442884 147486
rect 442644 147218 442646 147454
rect 442882 147218 442884 147454
rect 442644 147134 442884 147218
rect 442644 146898 442646 147134
rect 442882 146898 442884 147134
rect 442644 146866 442884 146898
rect 451644 147454 451884 147486
rect 451644 147218 451646 147454
rect 451882 147218 451884 147454
rect 451644 147134 451884 147218
rect 451644 146898 451646 147134
rect 451882 146898 451884 147134
rect 451644 146866 451884 146898
rect 460644 147454 460884 147486
rect 460644 147218 460646 147454
rect 460882 147218 460884 147454
rect 460644 147134 460884 147218
rect 460644 146898 460646 147134
rect 460882 146898 460884 147134
rect 460644 146866 460884 146898
rect 469644 147454 469884 147486
rect 469644 147218 469646 147454
rect 469882 147218 469884 147454
rect 469644 147134 469884 147218
rect 469644 146898 469646 147134
rect 469882 146898 469884 147134
rect 469644 146866 469884 146898
rect 471446 147454 471686 147486
rect 471446 147218 471448 147454
rect 471684 147218 471686 147454
rect 471446 147134 471686 147218
rect 471446 146898 471448 147134
rect 471684 146898 471686 147134
rect 471446 146866 471686 146898
rect 472818 147454 473058 147486
rect 472818 147218 472820 147454
rect 473056 147218 473058 147454
rect 472818 147134 473058 147218
rect 472818 146898 472820 147134
rect 473056 146898 473058 147134
rect 472818 146866 473058 146898
rect 473664 147454 473904 147486
rect 473664 147218 473666 147454
rect 473902 147218 473904 147454
rect 473664 147134 473904 147218
rect 473664 146898 473666 147134
rect 473902 146898 473904 147134
rect 473664 146866 473904 146898
rect 482664 147454 482904 147486
rect 482664 147218 482666 147454
rect 482902 147218 482904 147454
rect 482664 147134 482904 147218
rect 482664 146898 482666 147134
rect 482902 146898 482904 147134
rect 482664 146866 482904 146898
rect 491664 147454 491904 147486
rect 491664 147218 491666 147454
rect 491902 147218 491904 147454
rect 491664 147134 491904 147218
rect 491664 146898 491666 147134
rect 491902 146898 491904 147134
rect 491664 146866 491904 146898
rect 500664 147454 500904 147486
rect 500664 147218 500666 147454
rect 500902 147218 500904 147454
rect 500664 147134 500904 147218
rect 500664 146898 500666 147134
rect 500902 146898 500904 147134
rect 500664 146866 500904 146898
rect 509664 147454 509904 147486
rect 509664 147218 509666 147454
rect 509902 147218 509904 147454
rect 509664 147134 509904 147218
rect 509664 146898 509666 147134
rect 509902 146898 509904 147134
rect 509664 146866 509904 146898
rect 511466 147454 511706 147486
rect 511466 147218 511468 147454
rect 511704 147218 511706 147454
rect 511466 147134 511706 147218
rect 511466 146898 511468 147134
rect 511704 146898 511706 147134
rect 511466 146866 511706 146898
rect 512838 147454 513078 147486
rect 512838 147218 512840 147454
rect 513076 147218 513078 147454
rect 512838 147134 513078 147218
rect 512838 146898 512840 147134
rect 513076 146898 513078 147134
rect 512838 146866 513078 146898
rect 513684 147454 513924 147486
rect 513684 147218 513686 147454
rect 513922 147218 513924 147454
rect 513684 147134 513924 147218
rect 513684 146898 513686 147134
rect 513922 146898 513924 147134
rect 513684 146866 513924 146898
rect 522684 147454 522924 147486
rect 522684 147218 522686 147454
rect 522922 147218 522924 147454
rect 522684 147134 522924 147218
rect 522684 146898 522686 147134
rect 522922 146898 522924 147134
rect 522684 146866 522924 146898
rect 531684 147454 531924 147486
rect 531684 147218 531686 147454
rect 531922 147218 531924 147454
rect 531684 147134 531924 147218
rect 531684 146898 531686 147134
rect 531922 146898 531924 147134
rect 531684 146866 531924 146898
rect 540684 147454 540924 147486
rect 540684 147218 540686 147454
rect 540922 147218 540924 147454
rect 540684 147134 540924 147218
rect 540684 146898 540686 147134
rect 540922 146898 540924 147134
rect 540684 146866 540924 146898
rect 549684 147454 549924 147486
rect 549684 147218 549686 147454
rect 549922 147218 549924 147454
rect 549684 147134 549924 147218
rect 549684 146898 549686 147134
rect 549922 146898 549924 147134
rect 549684 146866 549924 146898
rect 551486 147454 551726 147486
rect 551486 147218 551488 147454
rect 551724 147218 551726 147454
rect 551486 147134 551726 147218
rect 551486 146898 551488 147134
rect 551724 146898 551726 147134
rect 551486 146866 551726 146898
rect 552858 147454 553098 147486
rect 552858 147218 552860 147454
rect 553096 147218 553098 147454
rect 552858 147134 553098 147218
rect 552858 146898 552860 147134
rect 553096 146898 553098 147134
rect 552858 146866 553098 146898
rect 553704 147454 553944 147486
rect 553704 147218 553706 147454
rect 553942 147218 553944 147454
rect 553704 147134 553944 147218
rect 553704 146898 553706 147134
rect 553942 146898 553944 147134
rect 553704 146866 553944 146898
rect 562704 147454 562944 147486
rect 562704 147218 562706 147454
rect 562942 147218 562944 147454
rect 562704 147134 562944 147218
rect 562704 146898 562706 147134
rect 562942 146898 562944 147134
rect 562704 146866 562944 146898
rect 571704 147454 571944 147486
rect 571704 147218 571706 147454
rect 571942 147218 571944 147454
rect 571704 147134 571944 147218
rect 571704 146898 571706 147134
rect 571942 146898 571944 147134
rect 571704 146866 571944 146898
rect 573474 147454 573714 147486
rect 573474 147218 573476 147454
rect 573712 147218 573714 147454
rect 573474 147134 573714 147218
rect 573474 146898 573476 147134
rect 573712 146898 573714 147134
rect 573474 146866 573714 146898
rect 578488 147454 579088 147486
rect 578488 147218 578670 147454
rect 578906 147218 579088 147454
rect 578488 147134 579088 147218
rect 578488 146898 578670 147134
rect 578906 146898 579088 147134
rect 578488 146866 579088 146898
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 4400 129454 5000 129486
rect 4400 129218 4582 129454
rect 4818 129218 5000 129454
rect 4400 129134 5000 129218
rect 4400 128898 4582 129134
rect 4818 128898 5000 129134
rect 4400 128866 5000 128898
rect 12230 129454 12470 129486
rect 12230 129218 12232 129454
rect 12468 129218 12470 129454
rect 12230 129134 12470 129218
rect 12230 128898 12232 129134
rect 12468 128898 12470 129134
rect 12230 128866 12470 128898
rect 13036 129454 13276 129486
rect 13036 129218 13038 129454
rect 13274 129218 13276 129454
rect 13036 129134 13276 129218
rect 13036 128898 13038 129134
rect 13274 128898 13276 129134
rect 13036 128866 13276 128898
rect 22036 129454 22276 129486
rect 22036 129218 22038 129454
rect 22274 129218 22276 129454
rect 22036 129134 22276 129218
rect 22036 128898 22038 129134
rect 22274 128898 22276 129134
rect 22036 128866 22276 128898
rect 27586 129454 27826 129486
rect 27586 129218 27588 129454
rect 27824 129218 27826 129454
rect 27586 129134 27826 129218
rect 27586 128898 27588 129134
rect 27824 128898 27826 129134
rect 27586 128866 27826 128898
rect 28238 129454 28478 129486
rect 28238 129218 28240 129454
rect 28476 129218 28478 129454
rect 28238 129134 28478 129218
rect 28238 128898 28240 129134
rect 28476 128898 28478 129134
rect 28238 128866 28478 128898
rect 29044 129454 29284 129486
rect 29044 129218 29046 129454
rect 29282 129218 29284 129454
rect 29044 129134 29284 129218
rect 29044 128898 29046 129134
rect 29282 128898 29284 129134
rect 29044 128866 29284 128898
rect 38044 129454 38284 129486
rect 38044 129218 38046 129454
rect 38282 129218 38284 129454
rect 38044 129134 38284 129218
rect 38044 128898 38046 129134
rect 38282 128898 38284 129134
rect 38044 128866 38284 128898
rect 47044 129454 47284 129486
rect 47044 129218 47046 129454
rect 47282 129218 47284 129454
rect 47044 129134 47284 129218
rect 47044 128898 47046 129134
rect 47282 128898 47284 129134
rect 47044 128866 47284 128898
rect 56044 129454 56284 129486
rect 56044 129218 56046 129454
rect 56282 129218 56284 129454
rect 56044 129134 56284 129218
rect 56044 128898 56046 129134
rect 56282 128898 56284 129134
rect 56044 128866 56284 128898
rect 65044 129454 65284 129486
rect 65044 129218 65046 129454
rect 65282 129218 65284 129454
rect 65044 129134 65284 129218
rect 65044 128898 65046 129134
rect 65282 128898 65284 129134
rect 65044 128866 65284 128898
rect 67606 129454 67846 129486
rect 67606 129218 67608 129454
rect 67844 129218 67846 129454
rect 67606 129134 67846 129218
rect 67606 128898 67608 129134
rect 67844 128898 67846 129134
rect 67606 128866 67846 128898
rect 68258 129454 68498 129486
rect 68258 129218 68260 129454
rect 68496 129218 68498 129454
rect 68258 129134 68498 129218
rect 68258 128898 68260 129134
rect 68496 128898 68498 129134
rect 68258 128866 68498 128898
rect 69064 129454 69304 129486
rect 69064 129218 69066 129454
rect 69302 129218 69304 129454
rect 69064 129134 69304 129218
rect 69064 128898 69066 129134
rect 69302 128898 69304 129134
rect 69064 128866 69304 128898
rect 78064 129454 78304 129486
rect 78064 129218 78066 129454
rect 78302 129218 78304 129454
rect 78064 129134 78304 129218
rect 78064 128898 78066 129134
rect 78302 128898 78304 129134
rect 78064 128866 78304 128898
rect 87064 129454 87304 129486
rect 87064 129218 87066 129454
rect 87302 129218 87304 129454
rect 87064 129134 87304 129218
rect 87064 128898 87066 129134
rect 87302 128898 87304 129134
rect 87064 128866 87304 128898
rect 96064 129454 96304 129486
rect 96064 129218 96066 129454
rect 96302 129218 96304 129454
rect 96064 129134 96304 129218
rect 96064 128898 96066 129134
rect 96302 128898 96304 129134
rect 96064 128866 96304 128898
rect 105064 129454 105304 129486
rect 105064 129218 105066 129454
rect 105302 129218 105304 129454
rect 105064 129134 105304 129218
rect 105064 128898 105066 129134
rect 105302 128898 105304 129134
rect 105064 128866 105304 128898
rect 107626 129454 107866 129486
rect 107626 129218 107628 129454
rect 107864 129218 107866 129454
rect 107626 129134 107866 129218
rect 107626 128898 107628 129134
rect 107864 128898 107866 129134
rect 107626 128866 107866 128898
rect 108278 129454 108518 129486
rect 108278 129218 108280 129454
rect 108516 129218 108518 129454
rect 108278 129134 108518 129218
rect 108278 128898 108280 129134
rect 108516 128898 108518 129134
rect 108278 128866 108518 128898
rect 109084 129454 109324 129486
rect 109084 129218 109086 129454
rect 109322 129218 109324 129454
rect 109084 129134 109324 129218
rect 109084 128898 109086 129134
rect 109322 128898 109324 129134
rect 109084 128866 109324 128898
rect 118084 129454 118324 129486
rect 118084 129218 118086 129454
rect 118322 129218 118324 129454
rect 118084 129134 118324 129218
rect 118084 128898 118086 129134
rect 118322 128898 118324 129134
rect 118084 128866 118324 128898
rect 127084 129454 127324 129486
rect 127084 129218 127086 129454
rect 127322 129218 127324 129454
rect 127084 129134 127324 129218
rect 127084 128898 127086 129134
rect 127322 128898 127324 129134
rect 127084 128866 127324 128898
rect 136084 129454 136324 129486
rect 136084 129218 136086 129454
rect 136322 129218 136324 129454
rect 136084 129134 136324 129218
rect 136084 128898 136086 129134
rect 136322 128898 136324 129134
rect 136084 128866 136324 128898
rect 145084 129454 145324 129486
rect 145084 129218 145086 129454
rect 145322 129218 145324 129454
rect 145084 129134 145324 129218
rect 145084 128898 145086 129134
rect 145322 128898 145324 129134
rect 145084 128866 145324 128898
rect 147646 129454 147886 129486
rect 147646 129218 147648 129454
rect 147884 129218 147886 129454
rect 147646 129134 147886 129218
rect 147646 128898 147648 129134
rect 147884 128898 147886 129134
rect 147646 128866 147886 128898
rect 149298 129454 149538 129486
rect 149298 129218 149300 129454
rect 149536 129218 149538 129454
rect 149298 129134 149538 129218
rect 149298 128898 149300 129134
rect 149536 128898 149538 129134
rect 149298 128866 149538 128898
rect 150104 129454 150344 129486
rect 150104 129218 150106 129454
rect 150342 129218 150344 129454
rect 150104 129134 150344 129218
rect 150104 128898 150106 129134
rect 150342 128898 150344 129134
rect 150104 128866 150344 128898
rect 159104 129454 159344 129486
rect 159104 129218 159106 129454
rect 159342 129218 159344 129454
rect 159104 129134 159344 129218
rect 159104 128898 159106 129134
rect 159342 128898 159344 129134
rect 159104 128866 159344 128898
rect 168104 129454 168344 129486
rect 168104 129218 168106 129454
rect 168342 129218 168344 129454
rect 168104 129134 168344 129218
rect 168104 128898 168106 129134
rect 168342 128898 168344 129134
rect 168104 128866 168344 128898
rect 177104 129454 177344 129486
rect 177104 129218 177106 129454
rect 177342 129218 177344 129454
rect 177104 129134 177344 129218
rect 177104 128898 177106 129134
rect 177342 128898 177344 129134
rect 177104 128866 177344 128898
rect 186104 129454 186344 129486
rect 186104 129218 186106 129454
rect 186342 129218 186344 129454
rect 186104 129134 186344 129218
rect 186104 128898 186106 129134
rect 186342 128898 186344 129134
rect 186104 128866 186344 128898
rect 188666 129454 188906 129486
rect 188666 129218 188668 129454
rect 188904 129218 188906 129454
rect 188666 129134 188906 129218
rect 188666 128898 188668 129134
rect 188904 128898 188906 129134
rect 188666 128866 188906 128898
rect 190318 129454 190558 129486
rect 190318 129218 190320 129454
rect 190556 129218 190558 129454
rect 190318 129134 190558 129218
rect 190318 128898 190320 129134
rect 190556 128898 190558 129134
rect 190318 128866 190558 128898
rect 191124 129454 191364 129486
rect 191124 129218 191126 129454
rect 191362 129218 191364 129454
rect 191124 129134 191364 129218
rect 191124 128898 191126 129134
rect 191362 128898 191364 129134
rect 191124 128866 191364 128898
rect 200124 129454 200364 129486
rect 200124 129218 200126 129454
rect 200362 129218 200364 129454
rect 200124 129134 200364 129218
rect 200124 128898 200126 129134
rect 200362 128898 200364 129134
rect 200124 128866 200364 128898
rect 209124 129454 209364 129486
rect 209124 129218 209126 129454
rect 209362 129218 209364 129454
rect 209124 129134 209364 129218
rect 209124 128898 209126 129134
rect 209362 128898 209364 129134
rect 209124 128866 209364 128898
rect 218124 129454 218364 129486
rect 218124 129218 218126 129454
rect 218362 129218 218364 129454
rect 218124 129134 218364 129218
rect 218124 128898 218126 129134
rect 218362 128898 218364 129134
rect 218124 128866 218364 128898
rect 227124 129454 227364 129486
rect 227124 129218 227126 129454
rect 227362 129218 227364 129454
rect 227124 129134 227364 129218
rect 227124 128898 227126 129134
rect 227362 128898 227364 129134
rect 227124 128866 227364 128898
rect 229686 129454 229926 129486
rect 229686 129218 229688 129454
rect 229924 129218 229926 129454
rect 229686 129134 229926 129218
rect 229686 128898 229688 129134
rect 229924 128898 229926 129134
rect 229686 128866 229926 128898
rect 230338 129454 230578 129486
rect 230338 129218 230340 129454
rect 230576 129218 230578 129454
rect 230338 129134 230578 129218
rect 230338 128898 230340 129134
rect 230576 128898 230578 129134
rect 230338 128866 230578 128898
rect 231144 129454 231384 129486
rect 231144 129218 231146 129454
rect 231382 129218 231384 129454
rect 231144 129134 231384 129218
rect 231144 128898 231146 129134
rect 231382 128898 231384 129134
rect 231144 128866 231384 128898
rect 240144 129454 240384 129486
rect 240144 129218 240146 129454
rect 240382 129218 240384 129454
rect 240144 129134 240384 129218
rect 240144 128898 240146 129134
rect 240382 128898 240384 129134
rect 240144 128866 240384 128898
rect 249144 129454 249384 129486
rect 249144 129218 249146 129454
rect 249382 129218 249384 129454
rect 249144 129134 249384 129218
rect 249144 128898 249146 129134
rect 249382 128898 249384 129134
rect 249144 128866 249384 128898
rect 258144 129454 258384 129486
rect 258144 129218 258146 129454
rect 258382 129218 258384 129454
rect 258144 129134 258384 129218
rect 258144 128898 258146 129134
rect 258382 128898 258384 129134
rect 258144 128866 258384 128898
rect 267144 129454 267384 129486
rect 267144 129218 267146 129454
rect 267382 129218 267384 129454
rect 267144 129134 267384 129218
rect 267144 128898 267146 129134
rect 267382 128898 267384 129134
rect 267144 128866 267384 128898
rect 269706 129454 269946 129486
rect 269706 129218 269708 129454
rect 269944 129218 269946 129454
rect 269706 129134 269946 129218
rect 269706 128898 269708 129134
rect 269944 128898 269946 129134
rect 269706 128866 269946 128898
rect 270358 129454 270598 129486
rect 270358 129218 270360 129454
rect 270596 129218 270598 129454
rect 270358 129134 270598 129218
rect 270358 128898 270360 129134
rect 270596 128898 270598 129134
rect 270358 128866 270598 128898
rect 271164 129454 271404 129486
rect 271164 129218 271166 129454
rect 271402 129218 271404 129454
rect 271164 129134 271404 129218
rect 271164 128898 271166 129134
rect 271402 128898 271404 129134
rect 271164 128866 271404 128898
rect 280164 129454 280404 129486
rect 280164 129218 280166 129454
rect 280402 129218 280404 129454
rect 280164 129134 280404 129218
rect 280164 128898 280166 129134
rect 280402 128898 280404 129134
rect 280164 128866 280404 128898
rect 289164 129454 289404 129486
rect 289164 129218 289166 129454
rect 289402 129218 289404 129454
rect 289164 129134 289404 129218
rect 289164 128898 289166 129134
rect 289402 128898 289404 129134
rect 289164 128866 289404 128898
rect 298164 129454 298404 129486
rect 298164 129218 298166 129454
rect 298402 129218 298404 129454
rect 298164 129134 298404 129218
rect 298164 128898 298166 129134
rect 298402 128898 298404 129134
rect 298164 128866 298404 128898
rect 307164 129454 307404 129486
rect 307164 129218 307166 129454
rect 307402 129218 307404 129454
rect 307164 129134 307404 129218
rect 307164 128898 307166 129134
rect 307402 128898 307404 129134
rect 307164 128866 307404 128898
rect 309726 129454 309966 129486
rect 309726 129218 309728 129454
rect 309964 129218 309966 129454
rect 309726 129134 309966 129218
rect 309726 128898 309728 129134
rect 309964 128898 309966 129134
rect 309726 128866 309966 128898
rect 311378 129454 311618 129486
rect 311378 129218 311380 129454
rect 311616 129218 311618 129454
rect 311378 129134 311618 129218
rect 311378 128898 311380 129134
rect 311616 128898 311618 129134
rect 311378 128866 311618 128898
rect 312184 129454 312424 129486
rect 312184 129218 312186 129454
rect 312422 129218 312424 129454
rect 312184 129134 312424 129218
rect 312184 128898 312186 129134
rect 312422 128898 312424 129134
rect 312184 128866 312424 128898
rect 321184 129454 321424 129486
rect 321184 129218 321186 129454
rect 321422 129218 321424 129454
rect 321184 129134 321424 129218
rect 321184 128898 321186 129134
rect 321422 128898 321424 129134
rect 321184 128866 321424 128898
rect 330184 129454 330424 129486
rect 330184 129218 330186 129454
rect 330422 129218 330424 129454
rect 330184 129134 330424 129218
rect 330184 128898 330186 129134
rect 330422 128898 330424 129134
rect 330184 128866 330424 128898
rect 339184 129454 339424 129486
rect 339184 129218 339186 129454
rect 339422 129218 339424 129454
rect 339184 129134 339424 129218
rect 339184 128898 339186 129134
rect 339422 128898 339424 129134
rect 339184 128866 339424 128898
rect 348184 129454 348424 129486
rect 348184 129218 348186 129454
rect 348422 129218 348424 129454
rect 348184 129134 348424 129218
rect 348184 128898 348186 129134
rect 348422 128898 348424 129134
rect 348184 128866 348424 128898
rect 350746 129454 350986 129486
rect 350746 129218 350748 129454
rect 350984 129218 350986 129454
rect 350746 129134 350986 129218
rect 350746 128898 350748 129134
rect 350984 128898 350986 129134
rect 350746 128866 350986 128898
rect 352398 129454 352638 129486
rect 352398 129218 352400 129454
rect 352636 129218 352638 129454
rect 352398 129134 352638 129218
rect 352398 128898 352400 129134
rect 352636 128898 352638 129134
rect 352398 128866 352638 128898
rect 353204 129454 353444 129486
rect 353204 129218 353206 129454
rect 353442 129218 353444 129454
rect 353204 129134 353444 129218
rect 353204 128898 353206 129134
rect 353442 128898 353444 129134
rect 353204 128866 353444 128898
rect 362204 129454 362444 129486
rect 362204 129218 362206 129454
rect 362442 129218 362444 129454
rect 362204 129134 362444 129218
rect 362204 128898 362206 129134
rect 362442 128898 362444 129134
rect 362204 128866 362444 128898
rect 371204 129454 371444 129486
rect 371204 129218 371206 129454
rect 371442 129218 371444 129454
rect 371204 129134 371444 129218
rect 371204 128898 371206 129134
rect 371442 128898 371444 129134
rect 371204 128866 371444 128898
rect 380204 129454 380444 129486
rect 380204 129218 380206 129454
rect 380442 129218 380444 129454
rect 380204 129134 380444 129218
rect 380204 128898 380206 129134
rect 380442 128898 380444 129134
rect 380204 128866 380444 128898
rect 389204 129454 389444 129486
rect 389204 129218 389206 129454
rect 389442 129218 389444 129454
rect 389204 129134 389444 129218
rect 389204 128898 389206 129134
rect 389442 128898 389444 129134
rect 389204 128866 389444 128898
rect 391766 129454 392006 129486
rect 391766 129218 391768 129454
rect 392004 129218 392006 129454
rect 391766 129134 392006 129218
rect 391766 128898 391768 129134
rect 392004 128898 392006 129134
rect 391766 128866 392006 128898
rect 392418 129454 392658 129486
rect 392418 129218 392420 129454
rect 392656 129218 392658 129454
rect 392418 129134 392658 129218
rect 392418 128898 392420 129134
rect 392656 128898 392658 129134
rect 392418 128866 392658 128898
rect 393224 129454 393464 129486
rect 393224 129218 393226 129454
rect 393462 129218 393464 129454
rect 393224 129134 393464 129218
rect 393224 128898 393226 129134
rect 393462 128898 393464 129134
rect 393224 128866 393464 128898
rect 402224 129454 402464 129486
rect 402224 129218 402226 129454
rect 402462 129218 402464 129454
rect 402224 129134 402464 129218
rect 402224 128898 402226 129134
rect 402462 128898 402464 129134
rect 402224 128866 402464 128898
rect 411224 129454 411464 129486
rect 411224 129218 411226 129454
rect 411462 129218 411464 129454
rect 411224 129134 411464 129218
rect 411224 128898 411226 129134
rect 411462 128898 411464 129134
rect 411224 128866 411464 128898
rect 420224 129454 420464 129486
rect 420224 129218 420226 129454
rect 420462 129218 420464 129454
rect 420224 129134 420464 129218
rect 420224 128898 420226 129134
rect 420462 128898 420464 129134
rect 420224 128866 420464 128898
rect 429224 129454 429464 129486
rect 429224 129218 429226 129454
rect 429462 129218 429464 129454
rect 429224 129134 429464 129218
rect 429224 128898 429226 129134
rect 429462 128898 429464 129134
rect 429224 128866 429464 128898
rect 431786 129454 432026 129486
rect 431786 129218 431788 129454
rect 432024 129218 432026 129454
rect 431786 129134 432026 129218
rect 431786 128898 431788 129134
rect 432024 128898 432026 129134
rect 431786 128866 432026 128898
rect 432438 129454 432678 129486
rect 432438 129218 432440 129454
rect 432676 129218 432678 129454
rect 432438 129134 432678 129218
rect 432438 128898 432440 129134
rect 432676 128898 432678 129134
rect 432438 128866 432678 128898
rect 433244 129454 433484 129486
rect 433244 129218 433246 129454
rect 433482 129218 433484 129454
rect 433244 129134 433484 129218
rect 433244 128898 433246 129134
rect 433482 128898 433484 129134
rect 433244 128866 433484 128898
rect 442244 129454 442484 129486
rect 442244 129218 442246 129454
rect 442482 129218 442484 129454
rect 442244 129134 442484 129218
rect 442244 128898 442246 129134
rect 442482 128898 442484 129134
rect 442244 128866 442484 128898
rect 451244 129454 451484 129486
rect 451244 129218 451246 129454
rect 451482 129218 451484 129454
rect 451244 129134 451484 129218
rect 451244 128898 451246 129134
rect 451482 128898 451484 129134
rect 451244 128866 451484 128898
rect 460244 129454 460484 129486
rect 460244 129218 460246 129454
rect 460482 129218 460484 129454
rect 460244 129134 460484 129218
rect 460244 128898 460246 129134
rect 460482 128898 460484 129134
rect 460244 128866 460484 128898
rect 469244 129454 469484 129486
rect 469244 129218 469246 129454
rect 469482 129218 469484 129454
rect 469244 129134 469484 129218
rect 469244 128898 469246 129134
rect 469482 128898 469484 129134
rect 469244 128866 469484 128898
rect 471806 129454 472046 129486
rect 471806 129218 471808 129454
rect 472044 129218 472046 129454
rect 471806 129134 472046 129218
rect 471806 128898 471808 129134
rect 472044 128898 472046 129134
rect 471806 128866 472046 128898
rect 472458 129454 472698 129486
rect 472458 129218 472460 129454
rect 472696 129218 472698 129454
rect 472458 129134 472698 129218
rect 472458 128898 472460 129134
rect 472696 128898 472698 129134
rect 472458 128866 472698 128898
rect 473264 129454 473504 129486
rect 473264 129218 473266 129454
rect 473502 129218 473504 129454
rect 473264 129134 473504 129218
rect 473264 128898 473266 129134
rect 473502 128898 473504 129134
rect 473264 128866 473504 128898
rect 482264 129454 482504 129486
rect 482264 129218 482266 129454
rect 482502 129218 482504 129454
rect 482264 129134 482504 129218
rect 482264 128898 482266 129134
rect 482502 128898 482504 129134
rect 482264 128866 482504 128898
rect 491264 129454 491504 129486
rect 491264 129218 491266 129454
rect 491502 129218 491504 129454
rect 491264 129134 491504 129218
rect 491264 128898 491266 129134
rect 491502 128898 491504 129134
rect 491264 128866 491504 128898
rect 500264 129454 500504 129486
rect 500264 129218 500266 129454
rect 500502 129218 500504 129454
rect 500264 129134 500504 129218
rect 500264 128898 500266 129134
rect 500502 128898 500504 129134
rect 500264 128866 500504 128898
rect 509264 129454 509504 129486
rect 509264 129218 509266 129454
rect 509502 129218 509504 129454
rect 509264 129134 509504 129218
rect 509264 128898 509266 129134
rect 509502 128898 509504 129134
rect 509264 128866 509504 128898
rect 511826 129454 512066 129486
rect 511826 129218 511828 129454
rect 512064 129218 512066 129454
rect 511826 129134 512066 129218
rect 511826 128898 511828 129134
rect 512064 128898 512066 129134
rect 511826 128866 512066 128898
rect 512478 129454 512718 129486
rect 512478 129218 512480 129454
rect 512716 129218 512718 129454
rect 512478 129134 512718 129218
rect 512478 128898 512480 129134
rect 512716 128898 512718 129134
rect 512478 128866 512718 128898
rect 513284 129454 513524 129486
rect 513284 129218 513286 129454
rect 513522 129218 513524 129454
rect 513284 129134 513524 129218
rect 513284 128898 513286 129134
rect 513522 128898 513524 129134
rect 513284 128866 513524 128898
rect 522284 129454 522524 129486
rect 522284 129218 522286 129454
rect 522522 129218 522524 129454
rect 522284 129134 522524 129218
rect 522284 128898 522286 129134
rect 522522 128898 522524 129134
rect 522284 128866 522524 128898
rect 531284 129454 531524 129486
rect 531284 129218 531286 129454
rect 531522 129218 531524 129454
rect 531284 129134 531524 129218
rect 531284 128898 531286 129134
rect 531522 128898 531524 129134
rect 531284 128866 531524 128898
rect 540284 129454 540524 129486
rect 540284 129218 540286 129454
rect 540522 129218 540524 129454
rect 540284 129134 540524 129218
rect 540284 128898 540286 129134
rect 540522 128898 540524 129134
rect 540284 128866 540524 128898
rect 549284 129454 549524 129486
rect 549284 129218 549286 129454
rect 549522 129218 549524 129454
rect 549284 129134 549524 129218
rect 549284 128898 549286 129134
rect 549522 128898 549524 129134
rect 549284 128866 549524 128898
rect 551846 129454 552086 129486
rect 551846 129218 551848 129454
rect 552084 129218 552086 129454
rect 551846 129134 552086 129218
rect 551846 128898 551848 129134
rect 552084 128898 552086 129134
rect 551846 128866 552086 128898
rect 552498 129454 552738 129486
rect 552498 129218 552500 129454
rect 552736 129218 552738 129454
rect 552498 129134 552738 129218
rect 552498 128898 552500 129134
rect 552736 128898 552738 129134
rect 552498 128866 552738 128898
rect 553304 129454 553544 129486
rect 553304 129218 553306 129454
rect 553542 129218 553544 129454
rect 553304 129134 553544 129218
rect 553304 128898 553306 129134
rect 553542 128898 553544 129134
rect 553304 128866 553544 128898
rect 562304 129454 562544 129486
rect 562304 129218 562306 129454
rect 562542 129218 562544 129454
rect 562304 129134 562544 129218
rect 562304 128898 562306 129134
rect 562542 128898 562544 129134
rect 562304 128866 562544 128898
rect 571304 129454 571544 129486
rect 571304 129218 571306 129454
rect 571542 129218 571544 129454
rect 571304 129134 571544 129218
rect 571304 128898 571306 129134
rect 571542 128898 571544 129134
rect 571304 128866 571544 128898
rect 573834 129454 574074 129486
rect 573834 129218 573836 129454
rect 574072 129218 574074 129454
rect 573834 129134 574074 129218
rect 573834 128898 573836 129134
rect 574072 128898 574074 129134
rect 573834 128866 574074 128898
rect 579288 129454 579888 129486
rect 579288 129218 579470 129454
rect 579706 129218 579888 129454
rect 579288 129134 579888 129218
rect 579288 128898 579470 129134
rect 579706 128898 579888 129134
rect 579288 128866 579888 128898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect 5200 111454 5800 111486
rect 5200 111218 5382 111454
rect 5618 111218 5800 111454
rect 5200 111134 5800 111218
rect 5200 110898 5382 111134
rect 5618 110898 5800 111134
rect 5200 110866 5800 110898
rect 12590 111454 12830 111486
rect 12590 111218 12592 111454
rect 12828 111218 12830 111454
rect 12590 111134 12830 111218
rect 12590 110898 12592 111134
rect 12828 110898 12830 111134
rect 12590 110866 12830 110898
rect 13436 111454 13676 111486
rect 13436 111218 13438 111454
rect 13674 111218 13676 111454
rect 13436 111134 13676 111218
rect 13436 110898 13438 111134
rect 13674 110898 13676 111134
rect 13436 110866 13676 110898
rect 22436 111454 22676 111486
rect 22436 111218 22438 111454
rect 22674 111218 22676 111454
rect 22436 111134 22676 111218
rect 22436 110898 22438 111134
rect 22674 110898 22676 111134
rect 22436 110866 22676 110898
rect 27226 111454 27466 111486
rect 27226 111218 27228 111454
rect 27464 111218 27466 111454
rect 27226 111134 27466 111218
rect 27226 110898 27228 111134
rect 27464 110898 27466 111134
rect 27226 110866 27466 110898
rect 28598 111454 28838 111486
rect 28598 111218 28600 111454
rect 28836 111218 28838 111454
rect 28598 111134 28838 111218
rect 28598 110898 28600 111134
rect 28836 110898 28838 111134
rect 28598 110866 28838 110898
rect 29444 111454 29684 111486
rect 29444 111218 29446 111454
rect 29682 111218 29684 111454
rect 29444 111134 29684 111218
rect 29444 110898 29446 111134
rect 29682 110898 29684 111134
rect 29444 110866 29684 110898
rect 38444 111454 38684 111486
rect 38444 111218 38446 111454
rect 38682 111218 38684 111454
rect 38444 111134 38684 111218
rect 38444 110898 38446 111134
rect 38682 110898 38684 111134
rect 38444 110866 38684 110898
rect 47444 111454 47684 111486
rect 47444 111218 47446 111454
rect 47682 111218 47684 111454
rect 47444 111134 47684 111218
rect 47444 110898 47446 111134
rect 47682 110898 47684 111134
rect 47444 110866 47684 110898
rect 56444 111454 56684 111486
rect 56444 111218 56446 111454
rect 56682 111218 56684 111454
rect 56444 111134 56684 111218
rect 56444 110898 56446 111134
rect 56682 110898 56684 111134
rect 56444 110866 56684 110898
rect 65444 111454 65684 111486
rect 65444 111218 65446 111454
rect 65682 111218 65684 111454
rect 65444 111134 65684 111218
rect 65444 110898 65446 111134
rect 65682 110898 65684 111134
rect 65444 110866 65684 110898
rect 67246 111454 67486 111486
rect 67246 111218 67248 111454
rect 67484 111218 67486 111454
rect 67246 111134 67486 111218
rect 67246 110898 67248 111134
rect 67484 110898 67486 111134
rect 67246 110866 67486 110898
rect 68618 111454 68858 111486
rect 68618 111218 68620 111454
rect 68856 111218 68858 111454
rect 68618 111134 68858 111218
rect 68618 110898 68620 111134
rect 68856 110898 68858 111134
rect 68618 110866 68858 110898
rect 69464 111454 69704 111486
rect 69464 111218 69466 111454
rect 69702 111218 69704 111454
rect 69464 111134 69704 111218
rect 69464 110898 69466 111134
rect 69702 110898 69704 111134
rect 69464 110866 69704 110898
rect 78464 111454 78704 111486
rect 78464 111218 78466 111454
rect 78702 111218 78704 111454
rect 78464 111134 78704 111218
rect 78464 110898 78466 111134
rect 78702 110898 78704 111134
rect 78464 110866 78704 110898
rect 87464 111454 87704 111486
rect 87464 111218 87466 111454
rect 87702 111218 87704 111454
rect 87464 111134 87704 111218
rect 87464 110898 87466 111134
rect 87702 110898 87704 111134
rect 87464 110866 87704 110898
rect 96464 111454 96704 111486
rect 96464 111218 96466 111454
rect 96702 111218 96704 111454
rect 96464 111134 96704 111218
rect 96464 110898 96466 111134
rect 96702 110898 96704 111134
rect 96464 110866 96704 110898
rect 105464 111454 105704 111486
rect 105464 111218 105466 111454
rect 105702 111218 105704 111454
rect 105464 111134 105704 111218
rect 105464 110898 105466 111134
rect 105702 110898 105704 111134
rect 105464 110866 105704 110898
rect 107266 111454 107506 111486
rect 107266 111218 107268 111454
rect 107504 111218 107506 111454
rect 107266 111134 107506 111218
rect 107266 110898 107268 111134
rect 107504 110898 107506 111134
rect 107266 110866 107506 110898
rect 108638 111454 108878 111486
rect 108638 111218 108640 111454
rect 108876 111218 108878 111454
rect 108638 111134 108878 111218
rect 108638 110898 108640 111134
rect 108876 110898 108878 111134
rect 108638 110866 108878 110898
rect 109484 111454 109724 111486
rect 109484 111218 109486 111454
rect 109722 111218 109724 111454
rect 109484 111134 109724 111218
rect 109484 110898 109486 111134
rect 109722 110898 109724 111134
rect 109484 110866 109724 110898
rect 118484 111454 118724 111486
rect 118484 111218 118486 111454
rect 118722 111218 118724 111454
rect 118484 111134 118724 111218
rect 118484 110898 118486 111134
rect 118722 110898 118724 111134
rect 118484 110866 118724 110898
rect 127484 111454 127724 111486
rect 127484 111218 127486 111454
rect 127722 111218 127724 111454
rect 127484 111134 127724 111218
rect 127484 110898 127486 111134
rect 127722 110898 127724 111134
rect 127484 110866 127724 110898
rect 136484 111454 136724 111486
rect 136484 111218 136486 111454
rect 136722 111218 136724 111454
rect 136484 111134 136724 111218
rect 136484 110898 136486 111134
rect 136722 110898 136724 111134
rect 136484 110866 136724 110898
rect 145484 111454 145724 111486
rect 145484 111218 145486 111454
rect 145722 111218 145724 111454
rect 145484 111134 145724 111218
rect 145484 110898 145486 111134
rect 145722 110898 145724 111134
rect 145484 110866 145724 110898
rect 147286 111454 147526 111486
rect 147286 111218 147288 111454
rect 147524 111218 147526 111454
rect 147286 111134 147526 111218
rect 147286 110898 147288 111134
rect 147524 110898 147526 111134
rect 147286 110866 147526 110898
rect 149658 111454 149898 111486
rect 149658 111218 149660 111454
rect 149896 111218 149898 111454
rect 149658 111134 149898 111218
rect 149658 110898 149660 111134
rect 149896 110898 149898 111134
rect 149658 110866 149898 110898
rect 150504 111454 150744 111486
rect 150504 111218 150506 111454
rect 150742 111218 150744 111454
rect 150504 111134 150744 111218
rect 150504 110898 150506 111134
rect 150742 110898 150744 111134
rect 150504 110866 150744 110898
rect 159504 111454 159744 111486
rect 159504 111218 159506 111454
rect 159742 111218 159744 111454
rect 159504 111134 159744 111218
rect 159504 110898 159506 111134
rect 159742 110898 159744 111134
rect 159504 110866 159744 110898
rect 168504 111454 168744 111486
rect 168504 111218 168506 111454
rect 168742 111218 168744 111454
rect 168504 111134 168744 111218
rect 168504 110898 168506 111134
rect 168742 110898 168744 111134
rect 168504 110866 168744 110898
rect 177504 111454 177744 111486
rect 177504 111218 177506 111454
rect 177742 111218 177744 111454
rect 177504 111134 177744 111218
rect 177504 110898 177506 111134
rect 177742 110898 177744 111134
rect 177504 110866 177744 110898
rect 186504 111454 186744 111486
rect 186504 111218 186506 111454
rect 186742 111218 186744 111454
rect 186504 111134 186744 111218
rect 186504 110898 186506 111134
rect 186742 110898 186744 111134
rect 186504 110866 186744 110898
rect 188306 111454 188546 111486
rect 188306 111218 188308 111454
rect 188544 111218 188546 111454
rect 188306 111134 188546 111218
rect 188306 110898 188308 111134
rect 188544 110898 188546 111134
rect 188306 110866 188546 110898
rect 190678 111454 190918 111486
rect 190678 111218 190680 111454
rect 190916 111218 190918 111454
rect 190678 111134 190918 111218
rect 190678 110898 190680 111134
rect 190916 110898 190918 111134
rect 190678 110866 190918 110898
rect 191524 111454 191764 111486
rect 191524 111218 191526 111454
rect 191762 111218 191764 111454
rect 191524 111134 191764 111218
rect 191524 110898 191526 111134
rect 191762 110898 191764 111134
rect 191524 110866 191764 110898
rect 200524 111454 200764 111486
rect 200524 111218 200526 111454
rect 200762 111218 200764 111454
rect 200524 111134 200764 111218
rect 200524 110898 200526 111134
rect 200762 110898 200764 111134
rect 200524 110866 200764 110898
rect 209524 111454 209764 111486
rect 209524 111218 209526 111454
rect 209762 111218 209764 111454
rect 209524 111134 209764 111218
rect 209524 110898 209526 111134
rect 209762 110898 209764 111134
rect 209524 110866 209764 110898
rect 218524 111454 218764 111486
rect 218524 111218 218526 111454
rect 218762 111218 218764 111454
rect 218524 111134 218764 111218
rect 218524 110898 218526 111134
rect 218762 110898 218764 111134
rect 218524 110866 218764 110898
rect 227524 111454 227764 111486
rect 227524 111218 227526 111454
rect 227762 111218 227764 111454
rect 227524 111134 227764 111218
rect 227524 110898 227526 111134
rect 227762 110898 227764 111134
rect 227524 110866 227764 110898
rect 229326 111454 229566 111486
rect 229326 111218 229328 111454
rect 229564 111218 229566 111454
rect 229326 111134 229566 111218
rect 229326 110898 229328 111134
rect 229564 110898 229566 111134
rect 229326 110866 229566 110898
rect 230698 111454 230938 111486
rect 230698 111218 230700 111454
rect 230936 111218 230938 111454
rect 230698 111134 230938 111218
rect 230698 110898 230700 111134
rect 230936 110898 230938 111134
rect 230698 110866 230938 110898
rect 231544 111454 231784 111486
rect 231544 111218 231546 111454
rect 231782 111218 231784 111454
rect 231544 111134 231784 111218
rect 231544 110898 231546 111134
rect 231782 110898 231784 111134
rect 231544 110866 231784 110898
rect 240544 111454 240784 111486
rect 240544 111218 240546 111454
rect 240782 111218 240784 111454
rect 240544 111134 240784 111218
rect 240544 110898 240546 111134
rect 240782 110898 240784 111134
rect 240544 110866 240784 110898
rect 249544 111454 249784 111486
rect 249544 111218 249546 111454
rect 249782 111218 249784 111454
rect 249544 111134 249784 111218
rect 249544 110898 249546 111134
rect 249782 110898 249784 111134
rect 249544 110866 249784 110898
rect 258544 111454 258784 111486
rect 258544 111218 258546 111454
rect 258782 111218 258784 111454
rect 258544 111134 258784 111218
rect 258544 110898 258546 111134
rect 258782 110898 258784 111134
rect 258544 110866 258784 110898
rect 267544 111454 267784 111486
rect 267544 111218 267546 111454
rect 267782 111218 267784 111454
rect 267544 111134 267784 111218
rect 267544 110898 267546 111134
rect 267782 110898 267784 111134
rect 267544 110866 267784 110898
rect 269346 111454 269586 111486
rect 269346 111218 269348 111454
rect 269584 111218 269586 111454
rect 269346 111134 269586 111218
rect 269346 110898 269348 111134
rect 269584 110898 269586 111134
rect 269346 110866 269586 110898
rect 270718 111454 270958 111486
rect 270718 111218 270720 111454
rect 270956 111218 270958 111454
rect 270718 111134 270958 111218
rect 270718 110898 270720 111134
rect 270956 110898 270958 111134
rect 270718 110866 270958 110898
rect 271564 111454 271804 111486
rect 271564 111218 271566 111454
rect 271802 111218 271804 111454
rect 271564 111134 271804 111218
rect 271564 110898 271566 111134
rect 271802 110898 271804 111134
rect 271564 110866 271804 110898
rect 280564 111454 280804 111486
rect 280564 111218 280566 111454
rect 280802 111218 280804 111454
rect 280564 111134 280804 111218
rect 280564 110898 280566 111134
rect 280802 110898 280804 111134
rect 280564 110866 280804 110898
rect 289564 111454 289804 111486
rect 289564 111218 289566 111454
rect 289802 111218 289804 111454
rect 289564 111134 289804 111218
rect 289564 110898 289566 111134
rect 289802 110898 289804 111134
rect 289564 110866 289804 110898
rect 298564 111454 298804 111486
rect 298564 111218 298566 111454
rect 298802 111218 298804 111454
rect 298564 111134 298804 111218
rect 298564 110898 298566 111134
rect 298802 110898 298804 111134
rect 298564 110866 298804 110898
rect 307564 111454 307804 111486
rect 307564 111218 307566 111454
rect 307802 111218 307804 111454
rect 307564 111134 307804 111218
rect 307564 110898 307566 111134
rect 307802 110898 307804 111134
rect 307564 110866 307804 110898
rect 309366 111454 309606 111486
rect 309366 111218 309368 111454
rect 309604 111218 309606 111454
rect 309366 111134 309606 111218
rect 309366 110898 309368 111134
rect 309604 110898 309606 111134
rect 309366 110866 309606 110898
rect 311738 111454 311978 111486
rect 311738 111218 311740 111454
rect 311976 111218 311978 111454
rect 311738 111134 311978 111218
rect 311738 110898 311740 111134
rect 311976 110898 311978 111134
rect 311738 110866 311978 110898
rect 312584 111454 312824 111486
rect 312584 111218 312586 111454
rect 312822 111218 312824 111454
rect 312584 111134 312824 111218
rect 312584 110898 312586 111134
rect 312822 110898 312824 111134
rect 312584 110866 312824 110898
rect 321584 111454 321824 111486
rect 321584 111218 321586 111454
rect 321822 111218 321824 111454
rect 321584 111134 321824 111218
rect 321584 110898 321586 111134
rect 321822 110898 321824 111134
rect 321584 110866 321824 110898
rect 330584 111454 330824 111486
rect 330584 111218 330586 111454
rect 330822 111218 330824 111454
rect 330584 111134 330824 111218
rect 330584 110898 330586 111134
rect 330822 110898 330824 111134
rect 330584 110866 330824 110898
rect 339584 111454 339824 111486
rect 339584 111218 339586 111454
rect 339822 111218 339824 111454
rect 339584 111134 339824 111218
rect 339584 110898 339586 111134
rect 339822 110898 339824 111134
rect 339584 110866 339824 110898
rect 348584 111454 348824 111486
rect 348584 111218 348586 111454
rect 348822 111218 348824 111454
rect 348584 111134 348824 111218
rect 348584 110898 348586 111134
rect 348822 110898 348824 111134
rect 348584 110866 348824 110898
rect 350386 111454 350626 111486
rect 350386 111218 350388 111454
rect 350624 111218 350626 111454
rect 350386 111134 350626 111218
rect 350386 110898 350388 111134
rect 350624 110898 350626 111134
rect 350386 110866 350626 110898
rect 352758 111454 352998 111486
rect 352758 111218 352760 111454
rect 352996 111218 352998 111454
rect 352758 111134 352998 111218
rect 352758 110898 352760 111134
rect 352996 110898 352998 111134
rect 352758 110866 352998 110898
rect 353604 111454 353844 111486
rect 353604 111218 353606 111454
rect 353842 111218 353844 111454
rect 353604 111134 353844 111218
rect 353604 110898 353606 111134
rect 353842 110898 353844 111134
rect 353604 110866 353844 110898
rect 362604 111454 362844 111486
rect 362604 111218 362606 111454
rect 362842 111218 362844 111454
rect 362604 111134 362844 111218
rect 362604 110898 362606 111134
rect 362842 110898 362844 111134
rect 362604 110866 362844 110898
rect 371604 111454 371844 111486
rect 371604 111218 371606 111454
rect 371842 111218 371844 111454
rect 371604 111134 371844 111218
rect 371604 110898 371606 111134
rect 371842 110898 371844 111134
rect 371604 110866 371844 110898
rect 380604 111454 380844 111486
rect 380604 111218 380606 111454
rect 380842 111218 380844 111454
rect 380604 111134 380844 111218
rect 380604 110898 380606 111134
rect 380842 110898 380844 111134
rect 380604 110866 380844 110898
rect 389604 111454 389844 111486
rect 389604 111218 389606 111454
rect 389842 111218 389844 111454
rect 389604 111134 389844 111218
rect 389604 110898 389606 111134
rect 389842 110898 389844 111134
rect 389604 110866 389844 110898
rect 391406 111454 391646 111486
rect 391406 111218 391408 111454
rect 391644 111218 391646 111454
rect 391406 111134 391646 111218
rect 391406 110898 391408 111134
rect 391644 110898 391646 111134
rect 391406 110866 391646 110898
rect 392778 111454 393018 111486
rect 392778 111218 392780 111454
rect 393016 111218 393018 111454
rect 392778 111134 393018 111218
rect 392778 110898 392780 111134
rect 393016 110898 393018 111134
rect 392778 110866 393018 110898
rect 393624 111454 393864 111486
rect 393624 111218 393626 111454
rect 393862 111218 393864 111454
rect 393624 111134 393864 111218
rect 393624 110898 393626 111134
rect 393862 110898 393864 111134
rect 393624 110866 393864 110898
rect 402624 111454 402864 111486
rect 402624 111218 402626 111454
rect 402862 111218 402864 111454
rect 402624 111134 402864 111218
rect 402624 110898 402626 111134
rect 402862 110898 402864 111134
rect 402624 110866 402864 110898
rect 411624 111454 411864 111486
rect 411624 111218 411626 111454
rect 411862 111218 411864 111454
rect 411624 111134 411864 111218
rect 411624 110898 411626 111134
rect 411862 110898 411864 111134
rect 411624 110866 411864 110898
rect 420624 111454 420864 111486
rect 420624 111218 420626 111454
rect 420862 111218 420864 111454
rect 420624 111134 420864 111218
rect 420624 110898 420626 111134
rect 420862 110898 420864 111134
rect 420624 110866 420864 110898
rect 429624 111454 429864 111486
rect 429624 111218 429626 111454
rect 429862 111218 429864 111454
rect 429624 111134 429864 111218
rect 429624 110898 429626 111134
rect 429862 110898 429864 111134
rect 429624 110866 429864 110898
rect 431426 111454 431666 111486
rect 431426 111218 431428 111454
rect 431664 111218 431666 111454
rect 431426 111134 431666 111218
rect 431426 110898 431428 111134
rect 431664 110898 431666 111134
rect 431426 110866 431666 110898
rect 432798 111454 433038 111486
rect 432798 111218 432800 111454
rect 433036 111218 433038 111454
rect 432798 111134 433038 111218
rect 432798 110898 432800 111134
rect 433036 110898 433038 111134
rect 432798 110866 433038 110898
rect 433644 111454 433884 111486
rect 433644 111218 433646 111454
rect 433882 111218 433884 111454
rect 433644 111134 433884 111218
rect 433644 110898 433646 111134
rect 433882 110898 433884 111134
rect 433644 110866 433884 110898
rect 442644 111454 442884 111486
rect 442644 111218 442646 111454
rect 442882 111218 442884 111454
rect 442644 111134 442884 111218
rect 442644 110898 442646 111134
rect 442882 110898 442884 111134
rect 442644 110866 442884 110898
rect 451644 111454 451884 111486
rect 451644 111218 451646 111454
rect 451882 111218 451884 111454
rect 451644 111134 451884 111218
rect 451644 110898 451646 111134
rect 451882 110898 451884 111134
rect 451644 110866 451884 110898
rect 460644 111454 460884 111486
rect 460644 111218 460646 111454
rect 460882 111218 460884 111454
rect 460644 111134 460884 111218
rect 460644 110898 460646 111134
rect 460882 110898 460884 111134
rect 460644 110866 460884 110898
rect 469644 111454 469884 111486
rect 469644 111218 469646 111454
rect 469882 111218 469884 111454
rect 469644 111134 469884 111218
rect 469644 110898 469646 111134
rect 469882 110898 469884 111134
rect 469644 110866 469884 110898
rect 471446 111454 471686 111486
rect 471446 111218 471448 111454
rect 471684 111218 471686 111454
rect 471446 111134 471686 111218
rect 471446 110898 471448 111134
rect 471684 110898 471686 111134
rect 471446 110866 471686 110898
rect 472818 111454 473058 111486
rect 472818 111218 472820 111454
rect 473056 111218 473058 111454
rect 472818 111134 473058 111218
rect 472818 110898 472820 111134
rect 473056 110898 473058 111134
rect 472818 110866 473058 110898
rect 473664 111454 473904 111486
rect 473664 111218 473666 111454
rect 473902 111218 473904 111454
rect 473664 111134 473904 111218
rect 473664 110898 473666 111134
rect 473902 110898 473904 111134
rect 473664 110866 473904 110898
rect 482664 111454 482904 111486
rect 482664 111218 482666 111454
rect 482902 111218 482904 111454
rect 482664 111134 482904 111218
rect 482664 110898 482666 111134
rect 482902 110898 482904 111134
rect 482664 110866 482904 110898
rect 491664 111454 491904 111486
rect 491664 111218 491666 111454
rect 491902 111218 491904 111454
rect 491664 111134 491904 111218
rect 491664 110898 491666 111134
rect 491902 110898 491904 111134
rect 491664 110866 491904 110898
rect 500664 111454 500904 111486
rect 500664 111218 500666 111454
rect 500902 111218 500904 111454
rect 500664 111134 500904 111218
rect 500664 110898 500666 111134
rect 500902 110898 500904 111134
rect 500664 110866 500904 110898
rect 509664 111454 509904 111486
rect 509664 111218 509666 111454
rect 509902 111218 509904 111454
rect 509664 111134 509904 111218
rect 509664 110898 509666 111134
rect 509902 110898 509904 111134
rect 509664 110866 509904 110898
rect 511466 111454 511706 111486
rect 511466 111218 511468 111454
rect 511704 111218 511706 111454
rect 511466 111134 511706 111218
rect 511466 110898 511468 111134
rect 511704 110898 511706 111134
rect 511466 110866 511706 110898
rect 512838 111454 513078 111486
rect 512838 111218 512840 111454
rect 513076 111218 513078 111454
rect 512838 111134 513078 111218
rect 512838 110898 512840 111134
rect 513076 110898 513078 111134
rect 512838 110866 513078 110898
rect 513684 111454 513924 111486
rect 513684 111218 513686 111454
rect 513922 111218 513924 111454
rect 513684 111134 513924 111218
rect 513684 110898 513686 111134
rect 513922 110898 513924 111134
rect 513684 110866 513924 110898
rect 522684 111454 522924 111486
rect 522684 111218 522686 111454
rect 522922 111218 522924 111454
rect 522684 111134 522924 111218
rect 522684 110898 522686 111134
rect 522922 110898 522924 111134
rect 522684 110866 522924 110898
rect 531684 111454 531924 111486
rect 531684 111218 531686 111454
rect 531922 111218 531924 111454
rect 531684 111134 531924 111218
rect 531684 110898 531686 111134
rect 531922 110898 531924 111134
rect 531684 110866 531924 110898
rect 540684 111454 540924 111486
rect 540684 111218 540686 111454
rect 540922 111218 540924 111454
rect 540684 111134 540924 111218
rect 540684 110898 540686 111134
rect 540922 110898 540924 111134
rect 540684 110866 540924 110898
rect 549684 111454 549924 111486
rect 549684 111218 549686 111454
rect 549922 111218 549924 111454
rect 549684 111134 549924 111218
rect 549684 110898 549686 111134
rect 549922 110898 549924 111134
rect 549684 110866 549924 110898
rect 551486 111454 551726 111486
rect 551486 111218 551488 111454
rect 551724 111218 551726 111454
rect 551486 111134 551726 111218
rect 551486 110898 551488 111134
rect 551724 110898 551726 111134
rect 551486 110866 551726 110898
rect 552858 111454 553098 111486
rect 552858 111218 552860 111454
rect 553096 111218 553098 111454
rect 552858 111134 553098 111218
rect 552858 110898 552860 111134
rect 553096 110898 553098 111134
rect 552858 110866 553098 110898
rect 553704 111454 553944 111486
rect 553704 111218 553706 111454
rect 553942 111218 553944 111454
rect 553704 111134 553944 111218
rect 553704 110898 553706 111134
rect 553942 110898 553944 111134
rect 553704 110866 553944 110898
rect 562704 111454 562944 111486
rect 562704 111218 562706 111454
rect 562942 111218 562944 111454
rect 562704 111134 562944 111218
rect 562704 110898 562706 111134
rect 562942 110898 562944 111134
rect 562704 110866 562944 110898
rect 571704 111454 571944 111486
rect 571704 111218 571706 111454
rect 571942 111218 571944 111454
rect 571704 111134 571944 111218
rect 571704 110898 571706 111134
rect 571942 110898 571944 111134
rect 571704 110866 571944 110898
rect 573474 111454 573714 111486
rect 573474 111218 573476 111454
rect 573712 111218 573714 111454
rect 573474 111134 573714 111218
rect 573474 110898 573476 111134
rect 573712 110898 573714 111134
rect 573474 110866 573714 110898
rect 578488 111454 579088 111486
rect 578488 111218 578670 111454
rect 578906 111218 579088 111454
rect 578488 111134 579088 111218
rect 578488 110898 578670 111134
rect 578906 110898 579088 111134
rect 578488 110866 579088 110898
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 4400 93454 5000 93486
rect 4400 93218 4582 93454
rect 4818 93218 5000 93454
rect 4400 93134 5000 93218
rect 4400 92898 4582 93134
rect 4818 92898 5000 93134
rect 4400 92866 5000 92898
rect 12230 93454 12470 93486
rect 12230 93218 12232 93454
rect 12468 93218 12470 93454
rect 12230 93134 12470 93218
rect 12230 92898 12232 93134
rect 12468 92898 12470 93134
rect 12230 92866 12470 92898
rect 13036 93454 13276 93486
rect 13036 93218 13038 93454
rect 13274 93218 13276 93454
rect 13036 93134 13276 93218
rect 13036 92898 13038 93134
rect 13274 92898 13276 93134
rect 13036 92866 13276 92898
rect 22036 93454 22276 93486
rect 22036 93218 22038 93454
rect 22274 93218 22276 93454
rect 22036 93134 22276 93218
rect 22036 92898 22038 93134
rect 22274 92898 22276 93134
rect 22036 92866 22276 92898
rect 27586 93454 27826 93486
rect 27586 93218 27588 93454
rect 27824 93218 27826 93454
rect 27586 93134 27826 93218
rect 27586 92898 27588 93134
rect 27824 92898 27826 93134
rect 27586 92866 27826 92898
rect 28238 93454 28478 93486
rect 28238 93218 28240 93454
rect 28476 93218 28478 93454
rect 28238 93134 28478 93218
rect 28238 92898 28240 93134
rect 28476 92898 28478 93134
rect 28238 92866 28478 92898
rect 29044 93454 29284 93486
rect 29044 93218 29046 93454
rect 29282 93218 29284 93454
rect 29044 93134 29284 93218
rect 29044 92898 29046 93134
rect 29282 92898 29284 93134
rect 29044 92866 29284 92898
rect 38044 93454 38284 93486
rect 38044 93218 38046 93454
rect 38282 93218 38284 93454
rect 38044 93134 38284 93218
rect 38044 92898 38046 93134
rect 38282 92898 38284 93134
rect 38044 92866 38284 92898
rect 47044 93454 47284 93486
rect 47044 93218 47046 93454
rect 47282 93218 47284 93454
rect 47044 93134 47284 93218
rect 47044 92898 47046 93134
rect 47282 92898 47284 93134
rect 47044 92866 47284 92898
rect 56044 93454 56284 93486
rect 56044 93218 56046 93454
rect 56282 93218 56284 93454
rect 56044 93134 56284 93218
rect 56044 92898 56046 93134
rect 56282 92898 56284 93134
rect 56044 92866 56284 92898
rect 65044 93454 65284 93486
rect 65044 93218 65046 93454
rect 65282 93218 65284 93454
rect 65044 93134 65284 93218
rect 65044 92898 65046 93134
rect 65282 92898 65284 93134
rect 65044 92866 65284 92898
rect 67606 93454 67846 93486
rect 67606 93218 67608 93454
rect 67844 93218 67846 93454
rect 67606 93134 67846 93218
rect 67606 92898 67608 93134
rect 67844 92898 67846 93134
rect 67606 92866 67846 92898
rect 68258 93454 68498 93486
rect 68258 93218 68260 93454
rect 68496 93218 68498 93454
rect 68258 93134 68498 93218
rect 68258 92898 68260 93134
rect 68496 92898 68498 93134
rect 68258 92866 68498 92898
rect 69064 93454 69304 93486
rect 69064 93218 69066 93454
rect 69302 93218 69304 93454
rect 69064 93134 69304 93218
rect 69064 92898 69066 93134
rect 69302 92898 69304 93134
rect 69064 92866 69304 92898
rect 78064 93454 78304 93486
rect 78064 93218 78066 93454
rect 78302 93218 78304 93454
rect 78064 93134 78304 93218
rect 78064 92898 78066 93134
rect 78302 92898 78304 93134
rect 78064 92866 78304 92898
rect 87064 93454 87304 93486
rect 87064 93218 87066 93454
rect 87302 93218 87304 93454
rect 87064 93134 87304 93218
rect 87064 92898 87066 93134
rect 87302 92898 87304 93134
rect 87064 92866 87304 92898
rect 96064 93454 96304 93486
rect 96064 93218 96066 93454
rect 96302 93218 96304 93454
rect 96064 93134 96304 93218
rect 96064 92898 96066 93134
rect 96302 92898 96304 93134
rect 96064 92866 96304 92898
rect 105064 93454 105304 93486
rect 105064 93218 105066 93454
rect 105302 93218 105304 93454
rect 105064 93134 105304 93218
rect 105064 92898 105066 93134
rect 105302 92898 105304 93134
rect 105064 92866 105304 92898
rect 107626 93454 107866 93486
rect 107626 93218 107628 93454
rect 107864 93218 107866 93454
rect 107626 93134 107866 93218
rect 107626 92898 107628 93134
rect 107864 92898 107866 93134
rect 107626 92866 107866 92898
rect 108278 93454 108518 93486
rect 108278 93218 108280 93454
rect 108516 93218 108518 93454
rect 108278 93134 108518 93218
rect 108278 92898 108280 93134
rect 108516 92898 108518 93134
rect 108278 92866 108518 92898
rect 109084 93454 109324 93486
rect 109084 93218 109086 93454
rect 109322 93218 109324 93454
rect 109084 93134 109324 93218
rect 109084 92898 109086 93134
rect 109322 92898 109324 93134
rect 109084 92866 109324 92898
rect 118084 93454 118324 93486
rect 118084 93218 118086 93454
rect 118322 93218 118324 93454
rect 118084 93134 118324 93218
rect 118084 92898 118086 93134
rect 118322 92898 118324 93134
rect 118084 92866 118324 92898
rect 127084 93454 127324 93486
rect 127084 93218 127086 93454
rect 127322 93218 127324 93454
rect 127084 93134 127324 93218
rect 127084 92898 127086 93134
rect 127322 92898 127324 93134
rect 127084 92866 127324 92898
rect 136084 93454 136324 93486
rect 136084 93218 136086 93454
rect 136322 93218 136324 93454
rect 136084 93134 136324 93218
rect 136084 92898 136086 93134
rect 136322 92898 136324 93134
rect 136084 92866 136324 92898
rect 145084 93454 145324 93486
rect 145084 93218 145086 93454
rect 145322 93218 145324 93454
rect 145084 93134 145324 93218
rect 145084 92898 145086 93134
rect 145322 92898 145324 93134
rect 145084 92866 145324 92898
rect 147646 93454 147886 93486
rect 147646 93218 147648 93454
rect 147884 93218 147886 93454
rect 147646 93134 147886 93218
rect 147646 92898 147648 93134
rect 147884 92898 147886 93134
rect 147646 92866 147886 92898
rect 149298 93454 149538 93486
rect 149298 93218 149300 93454
rect 149536 93218 149538 93454
rect 149298 93134 149538 93218
rect 149298 92898 149300 93134
rect 149536 92898 149538 93134
rect 149298 92866 149538 92898
rect 150104 93454 150344 93486
rect 150104 93218 150106 93454
rect 150342 93218 150344 93454
rect 150104 93134 150344 93218
rect 150104 92898 150106 93134
rect 150342 92898 150344 93134
rect 150104 92866 150344 92898
rect 159104 93454 159344 93486
rect 159104 93218 159106 93454
rect 159342 93218 159344 93454
rect 159104 93134 159344 93218
rect 159104 92898 159106 93134
rect 159342 92898 159344 93134
rect 159104 92866 159344 92898
rect 168104 93454 168344 93486
rect 168104 93218 168106 93454
rect 168342 93218 168344 93454
rect 168104 93134 168344 93218
rect 168104 92898 168106 93134
rect 168342 92898 168344 93134
rect 168104 92866 168344 92898
rect 177104 93454 177344 93486
rect 177104 93218 177106 93454
rect 177342 93218 177344 93454
rect 177104 93134 177344 93218
rect 177104 92898 177106 93134
rect 177342 92898 177344 93134
rect 177104 92866 177344 92898
rect 186104 93454 186344 93486
rect 186104 93218 186106 93454
rect 186342 93218 186344 93454
rect 186104 93134 186344 93218
rect 186104 92898 186106 93134
rect 186342 92898 186344 93134
rect 186104 92866 186344 92898
rect 188666 93454 188906 93486
rect 188666 93218 188668 93454
rect 188904 93218 188906 93454
rect 188666 93134 188906 93218
rect 188666 92898 188668 93134
rect 188904 92898 188906 93134
rect 188666 92866 188906 92898
rect 190318 93454 190558 93486
rect 190318 93218 190320 93454
rect 190556 93218 190558 93454
rect 190318 93134 190558 93218
rect 190318 92898 190320 93134
rect 190556 92898 190558 93134
rect 190318 92866 190558 92898
rect 191124 93454 191364 93486
rect 191124 93218 191126 93454
rect 191362 93218 191364 93454
rect 191124 93134 191364 93218
rect 191124 92898 191126 93134
rect 191362 92898 191364 93134
rect 191124 92866 191364 92898
rect 200124 93454 200364 93486
rect 200124 93218 200126 93454
rect 200362 93218 200364 93454
rect 200124 93134 200364 93218
rect 200124 92898 200126 93134
rect 200362 92898 200364 93134
rect 200124 92866 200364 92898
rect 209124 93454 209364 93486
rect 209124 93218 209126 93454
rect 209362 93218 209364 93454
rect 209124 93134 209364 93218
rect 209124 92898 209126 93134
rect 209362 92898 209364 93134
rect 209124 92866 209364 92898
rect 218124 93454 218364 93486
rect 218124 93218 218126 93454
rect 218362 93218 218364 93454
rect 218124 93134 218364 93218
rect 218124 92898 218126 93134
rect 218362 92898 218364 93134
rect 218124 92866 218364 92898
rect 227124 93454 227364 93486
rect 227124 93218 227126 93454
rect 227362 93218 227364 93454
rect 227124 93134 227364 93218
rect 227124 92898 227126 93134
rect 227362 92898 227364 93134
rect 227124 92866 227364 92898
rect 229686 93454 229926 93486
rect 229686 93218 229688 93454
rect 229924 93218 229926 93454
rect 229686 93134 229926 93218
rect 229686 92898 229688 93134
rect 229924 92898 229926 93134
rect 229686 92866 229926 92898
rect 230338 93454 230578 93486
rect 230338 93218 230340 93454
rect 230576 93218 230578 93454
rect 230338 93134 230578 93218
rect 230338 92898 230340 93134
rect 230576 92898 230578 93134
rect 230338 92866 230578 92898
rect 231144 93454 231384 93486
rect 231144 93218 231146 93454
rect 231382 93218 231384 93454
rect 231144 93134 231384 93218
rect 231144 92898 231146 93134
rect 231382 92898 231384 93134
rect 231144 92866 231384 92898
rect 240144 93454 240384 93486
rect 240144 93218 240146 93454
rect 240382 93218 240384 93454
rect 240144 93134 240384 93218
rect 240144 92898 240146 93134
rect 240382 92898 240384 93134
rect 240144 92866 240384 92898
rect 249144 93454 249384 93486
rect 249144 93218 249146 93454
rect 249382 93218 249384 93454
rect 249144 93134 249384 93218
rect 249144 92898 249146 93134
rect 249382 92898 249384 93134
rect 249144 92866 249384 92898
rect 258144 93454 258384 93486
rect 258144 93218 258146 93454
rect 258382 93218 258384 93454
rect 258144 93134 258384 93218
rect 258144 92898 258146 93134
rect 258382 92898 258384 93134
rect 258144 92866 258384 92898
rect 267144 93454 267384 93486
rect 267144 93218 267146 93454
rect 267382 93218 267384 93454
rect 267144 93134 267384 93218
rect 267144 92898 267146 93134
rect 267382 92898 267384 93134
rect 267144 92866 267384 92898
rect 269706 93454 269946 93486
rect 269706 93218 269708 93454
rect 269944 93218 269946 93454
rect 269706 93134 269946 93218
rect 269706 92898 269708 93134
rect 269944 92898 269946 93134
rect 269706 92866 269946 92898
rect 270358 93454 270598 93486
rect 270358 93218 270360 93454
rect 270596 93218 270598 93454
rect 270358 93134 270598 93218
rect 270358 92898 270360 93134
rect 270596 92898 270598 93134
rect 270358 92866 270598 92898
rect 271164 93454 271404 93486
rect 271164 93218 271166 93454
rect 271402 93218 271404 93454
rect 271164 93134 271404 93218
rect 271164 92898 271166 93134
rect 271402 92898 271404 93134
rect 271164 92866 271404 92898
rect 280164 93454 280404 93486
rect 280164 93218 280166 93454
rect 280402 93218 280404 93454
rect 280164 93134 280404 93218
rect 280164 92898 280166 93134
rect 280402 92898 280404 93134
rect 280164 92866 280404 92898
rect 289164 93454 289404 93486
rect 289164 93218 289166 93454
rect 289402 93218 289404 93454
rect 289164 93134 289404 93218
rect 289164 92898 289166 93134
rect 289402 92898 289404 93134
rect 289164 92866 289404 92898
rect 298164 93454 298404 93486
rect 298164 93218 298166 93454
rect 298402 93218 298404 93454
rect 298164 93134 298404 93218
rect 298164 92898 298166 93134
rect 298402 92898 298404 93134
rect 298164 92866 298404 92898
rect 307164 93454 307404 93486
rect 307164 93218 307166 93454
rect 307402 93218 307404 93454
rect 307164 93134 307404 93218
rect 307164 92898 307166 93134
rect 307402 92898 307404 93134
rect 307164 92866 307404 92898
rect 309726 93454 309966 93486
rect 309726 93218 309728 93454
rect 309964 93218 309966 93454
rect 309726 93134 309966 93218
rect 309726 92898 309728 93134
rect 309964 92898 309966 93134
rect 309726 92866 309966 92898
rect 311378 93454 311618 93486
rect 311378 93218 311380 93454
rect 311616 93218 311618 93454
rect 311378 93134 311618 93218
rect 311378 92898 311380 93134
rect 311616 92898 311618 93134
rect 311378 92866 311618 92898
rect 312184 93454 312424 93486
rect 312184 93218 312186 93454
rect 312422 93218 312424 93454
rect 312184 93134 312424 93218
rect 312184 92898 312186 93134
rect 312422 92898 312424 93134
rect 312184 92866 312424 92898
rect 321184 93454 321424 93486
rect 321184 93218 321186 93454
rect 321422 93218 321424 93454
rect 321184 93134 321424 93218
rect 321184 92898 321186 93134
rect 321422 92898 321424 93134
rect 321184 92866 321424 92898
rect 330184 93454 330424 93486
rect 330184 93218 330186 93454
rect 330422 93218 330424 93454
rect 330184 93134 330424 93218
rect 330184 92898 330186 93134
rect 330422 92898 330424 93134
rect 330184 92866 330424 92898
rect 339184 93454 339424 93486
rect 339184 93218 339186 93454
rect 339422 93218 339424 93454
rect 339184 93134 339424 93218
rect 339184 92898 339186 93134
rect 339422 92898 339424 93134
rect 339184 92866 339424 92898
rect 348184 93454 348424 93486
rect 348184 93218 348186 93454
rect 348422 93218 348424 93454
rect 348184 93134 348424 93218
rect 348184 92898 348186 93134
rect 348422 92898 348424 93134
rect 348184 92866 348424 92898
rect 350746 93454 350986 93486
rect 350746 93218 350748 93454
rect 350984 93218 350986 93454
rect 350746 93134 350986 93218
rect 350746 92898 350748 93134
rect 350984 92898 350986 93134
rect 350746 92866 350986 92898
rect 352398 93454 352638 93486
rect 352398 93218 352400 93454
rect 352636 93218 352638 93454
rect 352398 93134 352638 93218
rect 352398 92898 352400 93134
rect 352636 92898 352638 93134
rect 352398 92866 352638 92898
rect 353204 93454 353444 93486
rect 353204 93218 353206 93454
rect 353442 93218 353444 93454
rect 353204 93134 353444 93218
rect 353204 92898 353206 93134
rect 353442 92898 353444 93134
rect 353204 92866 353444 92898
rect 362204 93454 362444 93486
rect 362204 93218 362206 93454
rect 362442 93218 362444 93454
rect 362204 93134 362444 93218
rect 362204 92898 362206 93134
rect 362442 92898 362444 93134
rect 362204 92866 362444 92898
rect 371204 93454 371444 93486
rect 371204 93218 371206 93454
rect 371442 93218 371444 93454
rect 371204 93134 371444 93218
rect 371204 92898 371206 93134
rect 371442 92898 371444 93134
rect 371204 92866 371444 92898
rect 380204 93454 380444 93486
rect 380204 93218 380206 93454
rect 380442 93218 380444 93454
rect 380204 93134 380444 93218
rect 380204 92898 380206 93134
rect 380442 92898 380444 93134
rect 380204 92866 380444 92898
rect 389204 93454 389444 93486
rect 389204 93218 389206 93454
rect 389442 93218 389444 93454
rect 389204 93134 389444 93218
rect 389204 92898 389206 93134
rect 389442 92898 389444 93134
rect 389204 92866 389444 92898
rect 391766 93454 392006 93486
rect 391766 93218 391768 93454
rect 392004 93218 392006 93454
rect 391766 93134 392006 93218
rect 391766 92898 391768 93134
rect 392004 92898 392006 93134
rect 391766 92866 392006 92898
rect 392418 93454 392658 93486
rect 392418 93218 392420 93454
rect 392656 93218 392658 93454
rect 392418 93134 392658 93218
rect 392418 92898 392420 93134
rect 392656 92898 392658 93134
rect 392418 92866 392658 92898
rect 393224 93454 393464 93486
rect 393224 93218 393226 93454
rect 393462 93218 393464 93454
rect 393224 93134 393464 93218
rect 393224 92898 393226 93134
rect 393462 92898 393464 93134
rect 393224 92866 393464 92898
rect 402224 93454 402464 93486
rect 402224 93218 402226 93454
rect 402462 93218 402464 93454
rect 402224 93134 402464 93218
rect 402224 92898 402226 93134
rect 402462 92898 402464 93134
rect 402224 92866 402464 92898
rect 411224 93454 411464 93486
rect 411224 93218 411226 93454
rect 411462 93218 411464 93454
rect 411224 93134 411464 93218
rect 411224 92898 411226 93134
rect 411462 92898 411464 93134
rect 411224 92866 411464 92898
rect 420224 93454 420464 93486
rect 420224 93218 420226 93454
rect 420462 93218 420464 93454
rect 420224 93134 420464 93218
rect 420224 92898 420226 93134
rect 420462 92898 420464 93134
rect 420224 92866 420464 92898
rect 429224 93454 429464 93486
rect 429224 93218 429226 93454
rect 429462 93218 429464 93454
rect 429224 93134 429464 93218
rect 429224 92898 429226 93134
rect 429462 92898 429464 93134
rect 429224 92866 429464 92898
rect 431786 93454 432026 93486
rect 431786 93218 431788 93454
rect 432024 93218 432026 93454
rect 431786 93134 432026 93218
rect 431786 92898 431788 93134
rect 432024 92898 432026 93134
rect 431786 92866 432026 92898
rect 432438 93454 432678 93486
rect 432438 93218 432440 93454
rect 432676 93218 432678 93454
rect 432438 93134 432678 93218
rect 432438 92898 432440 93134
rect 432676 92898 432678 93134
rect 432438 92866 432678 92898
rect 433244 93454 433484 93486
rect 433244 93218 433246 93454
rect 433482 93218 433484 93454
rect 433244 93134 433484 93218
rect 433244 92898 433246 93134
rect 433482 92898 433484 93134
rect 433244 92866 433484 92898
rect 442244 93454 442484 93486
rect 442244 93218 442246 93454
rect 442482 93218 442484 93454
rect 442244 93134 442484 93218
rect 442244 92898 442246 93134
rect 442482 92898 442484 93134
rect 442244 92866 442484 92898
rect 451244 93454 451484 93486
rect 451244 93218 451246 93454
rect 451482 93218 451484 93454
rect 451244 93134 451484 93218
rect 451244 92898 451246 93134
rect 451482 92898 451484 93134
rect 451244 92866 451484 92898
rect 460244 93454 460484 93486
rect 460244 93218 460246 93454
rect 460482 93218 460484 93454
rect 460244 93134 460484 93218
rect 460244 92898 460246 93134
rect 460482 92898 460484 93134
rect 460244 92866 460484 92898
rect 469244 93454 469484 93486
rect 469244 93218 469246 93454
rect 469482 93218 469484 93454
rect 469244 93134 469484 93218
rect 469244 92898 469246 93134
rect 469482 92898 469484 93134
rect 469244 92866 469484 92898
rect 471806 93454 472046 93486
rect 471806 93218 471808 93454
rect 472044 93218 472046 93454
rect 471806 93134 472046 93218
rect 471806 92898 471808 93134
rect 472044 92898 472046 93134
rect 471806 92866 472046 92898
rect 472458 93454 472698 93486
rect 472458 93218 472460 93454
rect 472696 93218 472698 93454
rect 472458 93134 472698 93218
rect 472458 92898 472460 93134
rect 472696 92898 472698 93134
rect 472458 92866 472698 92898
rect 473264 93454 473504 93486
rect 473264 93218 473266 93454
rect 473502 93218 473504 93454
rect 473264 93134 473504 93218
rect 473264 92898 473266 93134
rect 473502 92898 473504 93134
rect 473264 92866 473504 92898
rect 482264 93454 482504 93486
rect 482264 93218 482266 93454
rect 482502 93218 482504 93454
rect 482264 93134 482504 93218
rect 482264 92898 482266 93134
rect 482502 92898 482504 93134
rect 482264 92866 482504 92898
rect 491264 93454 491504 93486
rect 491264 93218 491266 93454
rect 491502 93218 491504 93454
rect 491264 93134 491504 93218
rect 491264 92898 491266 93134
rect 491502 92898 491504 93134
rect 491264 92866 491504 92898
rect 500264 93454 500504 93486
rect 500264 93218 500266 93454
rect 500502 93218 500504 93454
rect 500264 93134 500504 93218
rect 500264 92898 500266 93134
rect 500502 92898 500504 93134
rect 500264 92866 500504 92898
rect 509264 93454 509504 93486
rect 509264 93218 509266 93454
rect 509502 93218 509504 93454
rect 509264 93134 509504 93218
rect 509264 92898 509266 93134
rect 509502 92898 509504 93134
rect 509264 92866 509504 92898
rect 511826 93454 512066 93486
rect 511826 93218 511828 93454
rect 512064 93218 512066 93454
rect 511826 93134 512066 93218
rect 511826 92898 511828 93134
rect 512064 92898 512066 93134
rect 511826 92866 512066 92898
rect 512478 93454 512718 93486
rect 512478 93218 512480 93454
rect 512716 93218 512718 93454
rect 512478 93134 512718 93218
rect 512478 92898 512480 93134
rect 512716 92898 512718 93134
rect 512478 92866 512718 92898
rect 513284 93454 513524 93486
rect 513284 93218 513286 93454
rect 513522 93218 513524 93454
rect 513284 93134 513524 93218
rect 513284 92898 513286 93134
rect 513522 92898 513524 93134
rect 513284 92866 513524 92898
rect 522284 93454 522524 93486
rect 522284 93218 522286 93454
rect 522522 93218 522524 93454
rect 522284 93134 522524 93218
rect 522284 92898 522286 93134
rect 522522 92898 522524 93134
rect 522284 92866 522524 92898
rect 531284 93454 531524 93486
rect 531284 93218 531286 93454
rect 531522 93218 531524 93454
rect 531284 93134 531524 93218
rect 531284 92898 531286 93134
rect 531522 92898 531524 93134
rect 531284 92866 531524 92898
rect 540284 93454 540524 93486
rect 540284 93218 540286 93454
rect 540522 93218 540524 93454
rect 540284 93134 540524 93218
rect 540284 92898 540286 93134
rect 540522 92898 540524 93134
rect 540284 92866 540524 92898
rect 549284 93454 549524 93486
rect 549284 93218 549286 93454
rect 549522 93218 549524 93454
rect 549284 93134 549524 93218
rect 549284 92898 549286 93134
rect 549522 92898 549524 93134
rect 549284 92866 549524 92898
rect 551846 93454 552086 93486
rect 551846 93218 551848 93454
rect 552084 93218 552086 93454
rect 551846 93134 552086 93218
rect 551846 92898 551848 93134
rect 552084 92898 552086 93134
rect 551846 92866 552086 92898
rect 552498 93454 552738 93486
rect 552498 93218 552500 93454
rect 552736 93218 552738 93454
rect 552498 93134 552738 93218
rect 552498 92898 552500 93134
rect 552736 92898 552738 93134
rect 552498 92866 552738 92898
rect 553304 93454 553544 93486
rect 553304 93218 553306 93454
rect 553542 93218 553544 93454
rect 553304 93134 553544 93218
rect 553304 92898 553306 93134
rect 553542 92898 553544 93134
rect 553304 92866 553544 92898
rect 562304 93454 562544 93486
rect 562304 93218 562306 93454
rect 562542 93218 562544 93454
rect 562304 93134 562544 93218
rect 562304 92898 562306 93134
rect 562542 92898 562544 93134
rect 562304 92866 562544 92898
rect 571304 93454 571544 93486
rect 571304 93218 571306 93454
rect 571542 93218 571544 93454
rect 571304 93134 571544 93218
rect 571304 92898 571306 93134
rect 571542 92898 571544 93134
rect 571304 92866 571544 92898
rect 573834 93454 574074 93486
rect 573834 93218 573836 93454
rect 574072 93218 574074 93454
rect 573834 93134 574074 93218
rect 573834 92898 573836 93134
rect 574072 92898 574074 93134
rect 573834 92866 574074 92898
rect 579288 93454 579888 93486
rect 579288 93218 579470 93454
rect 579706 93218 579888 93454
rect 579288 93134 579888 93218
rect 579288 92898 579470 93134
rect 579706 92898 579888 93134
rect 579288 92866 579888 92898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect 5200 75454 5800 75486
rect 5200 75218 5382 75454
rect 5618 75218 5800 75454
rect 5200 75134 5800 75218
rect 5200 74898 5382 75134
rect 5618 74898 5800 75134
rect 5200 74866 5800 74898
rect 12590 75454 12830 75486
rect 12590 75218 12592 75454
rect 12828 75218 12830 75454
rect 12590 75134 12830 75218
rect 12590 74898 12592 75134
rect 12828 74898 12830 75134
rect 12590 74866 12830 74898
rect 13436 75454 13676 75486
rect 13436 75218 13438 75454
rect 13674 75218 13676 75454
rect 13436 75134 13676 75218
rect 13436 74898 13438 75134
rect 13674 74898 13676 75134
rect 13436 74866 13676 74898
rect 22436 75454 22676 75486
rect 22436 75218 22438 75454
rect 22674 75218 22676 75454
rect 22436 75134 22676 75218
rect 22436 74898 22438 75134
rect 22674 74898 22676 75134
rect 22436 74866 22676 74898
rect 27226 75454 27466 75486
rect 27226 75218 27228 75454
rect 27464 75218 27466 75454
rect 27226 75134 27466 75218
rect 27226 74898 27228 75134
rect 27464 74898 27466 75134
rect 27226 74866 27466 74898
rect 28598 75454 28838 75486
rect 28598 75218 28600 75454
rect 28836 75218 28838 75454
rect 28598 75134 28838 75218
rect 28598 74898 28600 75134
rect 28836 74898 28838 75134
rect 28598 74866 28838 74898
rect 29444 75454 29684 75486
rect 29444 75218 29446 75454
rect 29682 75218 29684 75454
rect 29444 75134 29684 75218
rect 29444 74898 29446 75134
rect 29682 74898 29684 75134
rect 29444 74866 29684 74898
rect 38444 75454 38684 75486
rect 38444 75218 38446 75454
rect 38682 75218 38684 75454
rect 38444 75134 38684 75218
rect 38444 74898 38446 75134
rect 38682 74898 38684 75134
rect 38444 74866 38684 74898
rect 47444 75454 47684 75486
rect 47444 75218 47446 75454
rect 47682 75218 47684 75454
rect 47444 75134 47684 75218
rect 47444 74898 47446 75134
rect 47682 74898 47684 75134
rect 47444 74866 47684 74898
rect 56444 75454 56684 75486
rect 56444 75218 56446 75454
rect 56682 75218 56684 75454
rect 56444 75134 56684 75218
rect 56444 74898 56446 75134
rect 56682 74898 56684 75134
rect 56444 74866 56684 74898
rect 65444 75454 65684 75486
rect 65444 75218 65446 75454
rect 65682 75218 65684 75454
rect 65444 75134 65684 75218
rect 65444 74898 65446 75134
rect 65682 74898 65684 75134
rect 65444 74866 65684 74898
rect 67246 75454 67486 75486
rect 67246 75218 67248 75454
rect 67484 75218 67486 75454
rect 67246 75134 67486 75218
rect 67246 74898 67248 75134
rect 67484 74898 67486 75134
rect 67246 74866 67486 74898
rect 68618 75454 68858 75486
rect 68618 75218 68620 75454
rect 68856 75218 68858 75454
rect 68618 75134 68858 75218
rect 68618 74898 68620 75134
rect 68856 74898 68858 75134
rect 68618 74866 68858 74898
rect 69464 75454 69704 75486
rect 69464 75218 69466 75454
rect 69702 75218 69704 75454
rect 69464 75134 69704 75218
rect 69464 74898 69466 75134
rect 69702 74898 69704 75134
rect 69464 74866 69704 74898
rect 78464 75454 78704 75486
rect 78464 75218 78466 75454
rect 78702 75218 78704 75454
rect 78464 75134 78704 75218
rect 78464 74898 78466 75134
rect 78702 74898 78704 75134
rect 78464 74866 78704 74898
rect 87464 75454 87704 75486
rect 87464 75218 87466 75454
rect 87702 75218 87704 75454
rect 87464 75134 87704 75218
rect 87464 74898 87466 75134
rect 87702 74898 87704 75134
rect 87464 74866 87704 74898
rect 96464 75454 96704 75486
rect 96464 75218 96466 75454
rect 96702 75218 96704 75454
rect 96464 75134 96704 75218
rect 96464 74898 96466 75134
rect 96702 74898 96704 75134
rect 96464 74866 96704 74898
rect 105464 75454 105704 75486
rect 105464 75218 105466 75454
rect 105702 75218 105704 75454
rect 105464 75134 105704 75218
rect 105464 74898 105466 75134
rect 105702 74898 105704 75134
rect 105464 74866 105704 74898
rect 107266 75454 107506 75486
rect 107266 75218 107268 75454
rect 107504 75218 107506 75454
rect 107266 75134 107506 75218
rect 107266 74898 107268 75134
rect 107504 74898 107506 75134
rect 107266 74866 107506 74898
rect 108638 75454 108878 75486
rect 108638 75218 108640 75454
rect 108876 75218 108878 75454
rect 108638 75134 108878 75218
rect 108638 74898 108640 75134
rect 108876 74898 108878 75134
rect 108638 74866 108878 74898
rect 109484 75454 109724 75486
rect 109484 75218 109486 75454
rect 109722 75218 109724 75454
rect 109484 75134 109724 75218
rect 109484 74898 109486 75134
rect 109722 74898 109724 75134
rect 109484 74866 109724 74898
rect 118484 75454 118724 75486
rect 118484 75218 118486 75454
rect 118722 75218 118724 75454
rect 118484 75134 118724 75218
rect 118484 74898 118486 75134
rect 118722 74898 118724 75134
rect 118484 74866 118724 74898
rect 127484 75454 127724 75486
rect 127484 75218 127486 75454
rect 127722 75218 127724 75454
rect 127484 75134 127724 75218
rect 127484 74898 127486 75134
rect 127722 74898 127724 75134
rect 127484 74866 127724 74898
rect 136484 75454 136724 75486
rect 136484 75218 136486 75454
rect 136722 75218 136724 75454
rect 136484 75134 136724 75218
rect 136484 74898 136486 75134
rect 136722 74898 136724 75134
rect 136484 74866 136724 74898
rect 145484 75454 145724 75486
rect 145484 75218 145486 75454
rect 145722 75218 145724 75454
rect 145484 75134 145724 75218
rect 145484 74898 145486 75134
rect 145722 74898 145724 75134
rect 145484 74866 145724 74898
rect 147286 75454 147526 75486
rect 147286 75218 147288 75454
rect 147524 75218 147526 75454
rect 147286 75134 147526 75218
rect 147286 74898 147288 75134
rect 147524 74898 147526 75134
rect 147286 74866 147526 74898
rect 149658 75454 149898 75486
rect 149658 75218 149660 75454
rect 149896 75218 149898 75454
rect 149658 75134 149898 75218
rect 149658 74898 149660 75134
rect 149896 74898 149898 75134
rect 149658 74866 149898 74898
rect 150504 75454 150744 75486
rect 150504 75218 150506 75454
rect 150742 75218 150744 75454
rect 150504 75134 150744 75218
rect 150504 74898 150506 75134
rect 150742 74898 150744 75134
rect 150504 74866 150744 74898
rect 159504 75454 159744 75486
rect 159504 75218 159506 75454
rect 159742 75218 159744 75454
rect 159504 75134 159744 75218
rect 159504 74898 159506 75134
rect 159742 74898 159744 75134
rect 159504 74866 159744 74898
rect 168504 75454 168744 75486
rect 168504 75218 168506 75454
rect 168742 75218 168744 75454
rect 168504 75134 168744 75218
rect 168504 74898 168506 75134
rect 168742 74898 168744 75134
rect 168504 74866 168744 74898
rect 177504 75454 177744 75486
rect 177504 75218 177506 75454
rect 177742 75218 177744 75454
rect 177504 75134 177744 75218
rect 177504 74898 177506 75134
rect 177742 74898 177744 75134
rect 177504 74866 177744 74898
rect 186504 75454 186744 75486
rect 186504 75218 186506 75454
rect 186742 75218 186744 75454
rect 186504 75134 186744 75218
rect 186504 74898 186506 75134
rect 186742 74898 186744 75134
rect 186504 74866 186744 74898
rect 188306 75454 188546 75486
rect 188306 75218 188308 75454
rect 188544 75218 188546 75454
rect 188306 75134 188546 75218
rect 188306 74898 188308 75134
rect 188544 74898 188546 75134
rect 188306 74866 188546 74898
rect 190678 75454 190918 75486
rect 190678 75218 190680 75454
rect 190916 75218 190918 75454
rect 190678 75134 190918 75218
rect 190678 74898 190680 75134
rect 190916 74898 190918 75134
rect 190678 74866 190918 74898
rect 191524 75454 191764 75486
rect 191524 75218 191526 75454
rect 191762 75218 191764 75454
rect 191524 75134 191764 75218
rect 191524 74898 191526 75134
rect 191762 74898 191764 75134
rect 191524 74866 191764 74898
rect 200524 75454 200764 75486
rect 200524 75218 200526 75454
rect 200762 75218 200764 75454
rect 200524 75134 200764 75218
rect 200524 74898 200526 75134
rect 200762 74898 200764 75134
rect 200524 74866 200764 74898
rect 209524 75454 209764 75486
rect 209524 75218 209526 75454
rect 209762 75218 209764 75454
rect 209524 75134 209764 75218
rect 209524 74898 209526 75134
rect 209762 74898 209764 75134
rect 209524 74866 209764 74898
rect 218524 75454 218764 75486
rect 218524 75218 218526 75454
rect 218762 75218 218764 75454
rect 218524 75134 218764 75218
rect 218524 74898 218526 75134
rect 218762 74898 218764 75134
rect 218524 74866 218764 74898
rect 227524 75454 227764 75486
rect 227524 75218 227526 75454
rect 227762 75218 227764 75454
rect 227524 75134 227764 75218
rect 227524 74898 227526 75134
rect 227762 74898 227764 75134
rect 227524 74866 227764 74898
rect 229326 75454 229566 75486
rect 229326 75218 229328 75454
rect 229564 75218 229566 75454
rect 229326 75134 229566 75218
rect 229326 74898 229328 75134
rect 229564 74898 229566 75134
rect 229326 74866 229566 74898
rect 230698 75454 230938 75486
rect 230698 75218 230700 75454
rect 230936 75218 230938 75454
rect 230698 75134 230938 75218
rect 230698 74898 230700 75134
rect 230936 74898 230938 75134
rect 230698 74866 230938 74898
rect 231544 75454 231784 75486
rect 231544 75218 231546 75454
rect 231782 75218 231784 75454
rect 231544 75134 231784 75218
rect 231544 74898 231546 75134
rect 231782 74898 231784 75134
rect 231544 74866 231784 74898
rect 240544 75454 240784 75486
rect 240544 75218 240546 75454
rect 240782 75218 240784 75454
rect 240544 75134 240784 75218
rect 240544 74898 240546 75134
rect 240782 74898 240784 75134
rect 240544 74866 240784 74898
rect 249544 75454 249784 75486
rect 249544 75218 249546 75454
rect 249782 75218 249784 75454
rect 249544 75134 249784 75218
rect 249544 74898 249546 75134
rect 249782 74898 249784 75134
rect 249544 74866 249784 74898
rect 258544 75454 258784 75486
rect 258544 75218 258546 75454
rect 258782 75218 258784 75454
rect 258544 75134 258784 75218
rect 258544 74898 258546 75134
rect 258782 74898 258784 75134
rect 258544 74866 258784 74898
rect 267544 75454 267784 75486
rect 267544 75218 267546 75454
rect 267782 75218 267784 75454
rect 267544 75134 267784 75218
rect 267544 74898 267546 75134
rect 267782 74898 267784 75134
rect 267544 74866 267784 74898
rect 269346 75454 269586 75486
rect 269346 75218 269348 75454
rect 269584 75218 269586 75454
rect 269346 75134 269586 75218
rect 269346 74898 269348 75134
rect 269584 74898 269586 75134
rect 269346 74866 269586 74898
rect 270718 75454 270958 75486
rect 270718 75218 270720 75454
rect 270956 75218 270958 75454
rect 270718 75134 270958 75218
rect 270718 74898 270720 75134
rect 270956 74898 270958 75134
rect 270718 74866 270958 74898
rect 271564 75454 271804 75486
rect 271564 75218 271566 75454
rect 271802 75218 271804 75454
rect 271564 75134 271804 75218
rect 271564 74898 271566 75134
rect 271802 74898 271804 75134
rect 271564 74866 271804 74898
rect 280564 75454 280804 75486
rect 280564 75218 280566 75454
rect 280802 75218 280804 75454
rect 280564 75134 280804 75218
rect 280564 74898 280566 75134
rect 280802 74898 280804 75134
rect 280564 74866 280804 74898
rect 289564 75454 289804 75486
rect 289564 75218 289566 75454
rect 289802 75218 289804 75454
rect 289564 75134 289804 75218
rect 289564 74898 289566 75134
rect 289802 74898 289804 75134
rect 289564 74866 289804 74898
rect 298564 75454 298804 75486
rect 298564 75218 298566 75454
rect 298802 75218 298804 75454
rect 298564 75134 298804 75218
rect 298564 74898 298566 75134
rect 298802 74898 298804 75134
rect 298564 74866 298804 74898
rect 307564 75454 307804 75486
rect 307564 75218 307566 75454
rect 307802 75218 307804 75454
rect 307564 75134 307804 75218
rect 307564 74898 307566 75134
rect 307802 74898 307804 75134
rect 307564 74866 307804 74898
rect 309366 75454 309606 75486
rect 309366 75218 309368 75454
rect 309604 75218 309606 75454
rect 309366 75134 309606 75218
rect 309366 74898 309368 75134
rect 309604 74898 309606 75134
rect 309366 74866 309606 74898
rect 311738 75454 311978 75486
rect 311738 75218 311740 75454
rect 311976 75218 311978 75454
rect 311738 75134 311978 75218
rect 311738 74898 311740 75134
rect 311976 74898 311978 75134
rect 311738 74866 311978 74898
rect 312584 75454 312824 75486
rect 312584 75218 312586 75454
rect 312822 75218 312824 75454
rect 312584 75134 312824 75218
rect 312584 74898 312586 75134
rect 312822 74898 312824 75134
rect 312584 74866 312824 74898
rect 321584 75454 321824 75486
rect 321584 75218 321586 75454
rect 321822 75218 321824 75454
rect 321584 75134 321824 75218
rect 321584 74898 321586 75134
rect 321822 74898 321824 75134
rect 321584 74866 321824 74898
rect 330584 75454 330824 75486
rect 330584 75218 330586 75454
rect 330822 75218 330824 75454
rect 330584 75134 330824 75218
rect 330584 74898 330586 75134
rect 330822 74898 330824 75134
rect 330584 74866 330824 74898
rect 339584 75454 339824 75486
rect 339584 75218 339586 75454
rect 339822 75218 339824 75454
rect 339584 75134 339824 75218
rect 339584 74898 339586 75134
rect 339822 74898 339824 75134
rect 339584 74866 339824 74898
rect 348584 75454 348824 75486
rect 348584 75218 348586 75454
rect 348822 75218 348824 75454
rect 348584 75134 348824 75218
rect 348584 74898 348586 75134
rect 348822 74898 348824 75134
rect 348584 74866 348824 74898
rect 350386 75454 350626 75486
rect 350386 75218 350388 75454
rect 350624 75218 350626 75454
rect 350386 75134 350626 75218
rect 350386 74898 350388 75134
rect 350624 74898 350626 75134
rect 350386 74866 350626 74898
rect 352758 75454 352998 75486
rect 352758 75218 352760 75454
rect 352996 75218 352998 75454
rect 352758 75134 352998 75218
rect 352758 74898 352760 75134
rect 352996 74898 352998 75134
rect 352758 74866 352998 74898
rect 353604 75454 353844 75486
rect 353604 75218 353606 75454
rect 353842 75218 353844 75454
rect 353604 75134 353844 75218
rect 353604 74898 353606 75134
rect 353842 74898 353844 75134
rect 353604 74866 353844 74898
rect 362604 75454 362844 75486
rect 362604 75218 362606 75454
rect 362842 75218 362844 75454
rect 362604 75134 362844 75218
rect 362604 74898 362606 75134
rect 362842 74898 362844 75134
rect 362604 74866 362844 74898
rect 371604 75454 371844 75486
rect 371604 75218 371606 75454
rect 371842 75218 371844 75454
rect 371604 75134 371844 75218
rect 371604 74898 371606 75134
rect 371842 74898 371844 75134
rect 371604 74866 371844 74898
rect 380604 75454 380844 75486
rect 380604 75218 380606 75454
rect 380842 75218 380844 75454
rect 380604 75134 380844 75218
rect 380604 74898 380606 75134
rect 380842 74898 380844 75134
rect 380604 74866 380844 74898
rect 389604 75454 389844 75486
rect 389604 75218 389606 75454
rect 389842 75218 389844 75454
rect 389604 75134 389844 75218
rect 389604 74898 389606 75134
rect 389842 74898 389844 75134
rect 389604 74866 389844 74898
rect 391406 75454 391646 75486
rect 391406 75218 391408 75454
rect 391644 75218 391646 75454
rect 391406 75134 391646 75218
rect 391406 74898 391408 75134
rect 391644 74898 391646 75134
rect 391406 74866 391646 74898
rect 392778 75454 393018 75486
rect 392778 75218 392780 75454
rect 393016 75218 393018 75454
rect 392778 75134 393018 75218
rect 392778 74898 392780 75134
rect 393016 74898 393018 75134
rect 392778 74866 393018 74898
rect 393624 75454 393864 75486
rect 393624 75218 393626 75454
rect 393862 75218 393864 75454
rect 393624 75134 393864 75218
rect 393624 74898 393626 75134
rect 393862 74898 393864 75134
rect 393624 74866 393864 74898
rect 402624 75454 402864 75486
rect 402624 75218 402626 75454
rect 402862 75218 402864 75454
rect 402624 75134 402864 75218
rect 402624 74898 402626 75134
rect 402862 74898 402864 75134
rect 402624 74866 402864 74898
rect 411624 75454 411864 75486
rect 411624 75218 411626 75454
rect 411862 75218 411864 75454
rect 411624 75134 411864 75218
rect 411624 74898 411626 75134
rect 411862 74898 411864 75134
rect 411624 74866 411864 74898
rect 420624 75454 420864 75486
rect 420624 75218 420626 75454
rect 420862 75218 420864 75454
rect 420624 75134 420864 75218
rect 420624 74898 420626 75134
rect 420862 74898 420864 75134
rect 420624 74866 420864 74898
rect 429624 75454 429864 75486
rect 429624 75218 429626 75454
rect 429862 75218 429864 75454
rect 429624 75134 429864 75218
rect 429624 74898 429626 75134
rect 429862 74898 429864 75134
rect 429624 74866 429864 74898
rect 431426 75454 431666 75486
rect 431426 75218 431428 75454
rect 431664 75218 431666 75454
rect 431426 75134 431666 75218
rect 431426 74898 431428 75134
rect 431664 74898 431666 75134
rect 431426 74866 431666 74898
rect 432798 75454 433038 75486
rect 432798 75218 432800 75454
rect 433036 75218 433038 75454
rect 432798 75134 433038 75218
rect 432798 74898 432800 75134
rect 433036 74898 433038 75134
rect 432798 74866 433038 74898
rect 433644 75454 433884 75486
rect 433644 75218 433646 75454
rect 433882 75218 433884 75454
rect 433644 75134 433884 75218
rect 433644 74898 433646 75134
rect 433882 74898 433884 75134
rect 433644 74866 433884 74898
rect 442644 75454 442884 75486
rect 442644 75218 442646 75454
rect 442882 75218 442884 75454
rect 442644 75134 442884 75218
rect 442644 74898 442646 75134
rect 442882 74898 442884 75134
rect 442644 74866 442884 74898
rect 451644 75454 451884 75486
rect 451644 75218 451646 75454
rect 451882 75218 451884 75454
rect 451644 75134 451884 75218
rect 451644 74898 451646 75134
rect 451882 74898 451884 75134
rect 451644 74866 451884 74898
rect 460644 75454 460884 75486
rect 460644 75218 460646 75454
rect 460882 75218 460884 75454
rect 460644 75134 460884 75218
rect 460644 74898 460646 75134
rect 460882 74898 460884 75134
rect 460644 74866 460884 74898
rect 469644 75454 469884 75486
rect 469644 75218 469646 75454
rect 469882 75218 469884 75454
rect 469644 75134 469884 75218
rect 469644 74898 469646 75134
rect 469882 74898 469884 75134
rect 469644 74866 469884 74898
rect 471446 75454 471686 75486
rect 471446 75218 471448 75454
rect 471684 75218 471686 75454
rect 471446 75134 471686 75218
rect 471446 74898 471448 75134
rect 471684 74898 471686 75134
rect 471446 74866 471686 74898
rect 472818 75454 473058 75486
rect 472818 75218 472820 75454
rect 473056 75218 473058 75454
rect 472818 75134 473058 75218
rect 472818 74898 472820 75134
rect 473056 74898 473058 75134
rect 472818 74866 473058 74898
rect 473664 75454 473904 75486
rect 473664 75218 473666 75454
rect 473902 75218 473904 75454
rect 473664 75134 473904 75218
rect 473664 74898 473666 75134
rect 473902 74898 473904 75134
rect 473664 74866 473904 74898
rect 482664 75454 482904 75486
rect 482664 75218 482666 75454
rect 482902 75218 482904 75454
rect 482664 75134 482904 75218
rect 482664 74898 482666 75134
rect 482902 74898 482904 75134
rect 482664 74866 482904 74898
rect 491664 75454 491904 75486
rect 491664 75218 491666 75454
rect 491902 75218 491904 75454
rect 491664 75134 491904 75218
rect 491664 74898 491666 75134
rect 491902 74898 491904 75134
rect 491664 74866 491904 74898
rect 500664 75454 500904 75486
rect 500664 75218 500666 75454
rect 500902 75218 500904 75454
rect 500664 75134 500904 75218
rect 500664 74898 500666 75134
rect 500902 74898 500904 75134
rect 500664 74866 500904 74898
rect 509664 75454 509904 75486
rect 509664 75218 509666 75454
rect 509902 75218 509904 75454
rect 509664 75134 509904 75218
rect 509664 74898 509666 75134
rect 509902 74898 509904 75134
rect 509664 74866 509904 74898
rect 511466 75454 511706 75486
rect 511466 75218 511468 75454
rect 511704 75218 511706 75454
rect 511466 75134 511706 75218
rect 511466 74898 511468 75134
rect 511704 74898 511706 75134
rect 511466 74866 511706 74898
rect 512838 75454 513078 75486
rect 512838 75218 512840 75454
rect 513076 75218 513078 75454
rect 512838 75134 513078 75218
rect 512838 74898 512840 75134
rect 513076 74898 513078 75134
rect 512838 74866 513078 74898
rect 513684 75454 513924 75486
rect 513684 75218 513686 75454
rect 513922 75218 513924 75454
rect 513684 75134 513924 75218
rect 513684 74898 513686 75134
rect 513922 74898 513924 75134
rect 513684 74866 513924 74898
rect 522684 75454 522924 75486
rect 522684 75218 522686 75454
rect 522922 75218 522924 75454
rect 522684 75134 522924 75218
rect 522684 74898 522686 75134
rect 522922 74898 522924 75134
rect 522684 74866 522924 74898
rect 531684 75454 531924 75486
rect 531684 75218 531686 75454
rect 531922 75218 531924 75454
rect 531684 75134 531924 75218
rect 531684 74898 531686 75134
rect 531922 74898 531924 75134
rect 531684 74866 531924 74898
rect 540684 75454 540924 75486
rect 540684 75218 540686 75454
rect 540922 75218 540924 75454
rect 540684 75134 540924 75218
rect 540684 74898 540686 75134
rect 540922 74898 540924 75134
rect 540684 74866 540924 74898
rect 549684 75454 549924 75486
rect 549684 75218 549686 75454
rect 549922 75218 549924 75454
rect 549684 75134 549924 75218
rect 549684 74898 549686 75134
rect 549922 74898 549924 75134
rect 549684 74866 549924 74898
rect 551486 75454 551726 75486
rect 551486 75218 551488 75454
rect 551724 75218 551726 75454
rect 551486 75134 551726 75218
rect 551486 74898 551488 75134
rect 551724 74898 551726 75134
rect 551486 74866 551726 74898
rect 552858 75454 553098 75486
rect 552858 75218 552860 75454
rect 553096 75218 553098 75454
rect 552858 75134 553098 75218
rect 552858 74898 552860 75134
rect 553096 74898 553098 75134
rect 552858 74866 553098 74898
rect 553704 75454 553944 75486
rect 553704 75218 553706 75454
rect 553942 75218 553944 75454
rect 553704 75134 553944 75218
rect 553704 74898 553706 75134
rect 553942 74898 553944 75134
rect 553704 74866 553944 74898
rect 562704 75454 562944 75486
rect 562704 75218 562706 75454
rect 562942 75218 562944 75454
rect 562704 75134 562944 75218
rect 562704 74898 562706 75134
rect 562942 74898 562944 75134
rect 562704 74866 562944 74898
rect 571704 75454 571944 75486
rect 571704 75218 571706 75454
rect 571942 75218 571944 75454
rect 571704 75134 571944 75218
rect 571704 74898 571706 75134
rect 571942 74898 571944 75134
rect 571704 74866 571944 74898
rect 573474 75454 573714 75486
rect 573474 75218 573476 75454
rect 573712 75218 573714 75454
rect 573474 75134 573714 75218
rect 573474 74898 573476 75134
rect 573712 74898 573714 75134
rect 573474 74866 573714 74898
rect 578488 75454 579088 75486
rect 578488 75218 578670 75454
rect 578906 75218 579088 75454
rect 578488 75134 579088 75218
rect 578488 74898 578670 75134
rect 578906 74898 579088 75134
rect 578488 74866 579088 74898
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 4400 57454 5000 57486
rect 4400 57218 4582 57454
rect 4818 57218 5000 57454
rect 4400 57134 5000 57218
rect 4400 56898 4582 57134
rect 4818 56898 5000 57134
rect 4400 56866 5000 56898
rect 28238 57454 28478 57486
rect 28238 57218 28240 57454
rect 28476 57218 28478 57454
rect 28238 57134 28478 57218
rect 28238 56898 28240 57134
rect 28476 56898 28478 57134
rect 28238 56866 28478 56898
rect 29044 57454 29284 57486
rect 29044 57218 29046 57454
rect 29282 57218 29284 57454
rect 29044 57134 29284 57218
rect 29044 56898 29046 57134
rect 29282 56898 29284 57134
rect 29044 56866 29284 56898
rect 38044 57454 38284 57486
rect 38044 57218 38046 57454
rect 38282 57218 38284 57454
rect 38044 57134 38284 57218
rect 38044 56898 38046 57134
rect 38282 56898 38284 57134
rect 38044 56866 38284 56898
rect 47044 57454 47284 57486
rect 47044 57218 47046 57454
rect 47282 57218 47284 57454
rect 47044 57134 47284 57218
rect 47044 56898 47046 57134
rect 47282 56898 47284 57134
rect 47044 56866 47284 56898
rect 56044 57454 56284 57486
rect 56044 57218 56046 57454
rect 56282 57218 56284 57454
rect 56044 57134 56284 57218
rect 56044 56898 56046 57134
rect 56282 56898 56284 57134
rect 56044 56866 56284 56898
rect 65044 57454 65284 57486
rect 65044 57218 65046 57454
rect 65282 57218 65284 57454
rect 65044 57134 65284 57218
rect 65044 56898 65046 57134
rect 65282 56898 65284 57134
rect 65044 56866 65284 56898
rect 67606 57454 67846 57486
rect 67606 57218 67608 57454
rect 67844 57218 67846 57454
rect 67606 57134 67846 57218
rect 67606 56898 67608 57134
rect 67844 56898 67846 57134
rect 67606 56866 67846 56898
rect 68258 57454 68498 57486
rect 68258 57218 68260 57454
rect 68496 57218 68498 57454
rect 68258 57134 68498 57218
rect 68258 56898 68260 57134
rect 68496 56898 68498 57134
rect 68258 56866 68498 56898
rect 69064 57454 69304 57486
rect 69064 57218 69066 57454
rect 69302 57218 69304 57454
rect 69064 57134 69304 57218
rect 69064 56898 69066 57134
rect 69302 56898 69304 57134
rect 69064 56866 69304 56898
rect 78064 57454 78304 57486
rect 78064 57218 78066 57454
rect 78302 57218 78304 57454
rect 78064 57134 78304 57218
rect 78064 56898 78066 57134
rect 78302 56898 78304 57134
rect 78064 56866 78304 56898
rect 87064 57454 87304 57486
rect 87064 57218 87066 57454
rect 87302 57218 87304 57454
rect 87064 57134 87304 57218
rect 87064 56898 87066 57134
rect 87302 56898 87304 57134
rect 87064 56866 87304 56898
rect 96064 57454 96304 57486
rect 96064 57218 96066 57454
rect 96302 57218 96304 57454
rect 96064 57134 96304 57218
rect 96064 56898 96066 57134
rect 96302 56898 96304 57134
rect 96064 56866 96304 56898
rect 105064 57454 105304 57486
rect 105064 57218 105066 57454
rect 105302 57218 105304 57454
rect 105064 57134 105304 57218
rect 105064 56898 105066 57134
rect 105302 56898 105304 57134
rect 105064 56866 105304 56898
rect 107626 57454 107866 57486
rect 107626 57218 107628 57454
rect 107864 57218 107866 57454
rect 107626 57134 107866 57218
rect 107626 56898 107628 57134
rect 107864 56898 107866 57134
rect 107626 56866 107866 56898
rect 108278 57454 108518 57486
rect 108278 57218 108280 57454
rect 108516 57218 108518 57454
rect 108278 57134 108518 57218
rect 108278 56898 108280 57134
rect 108516 56898 108518 57134
rect 108278 56866 108518 56898
rect 109084 57454 109324 57486
rect 109084 57218 109086 57454
rect 109322 57218 109324 57454
rect 109084 57134 109324 57218
rect 109084 56898 109086 57134
rect 109322 56898 109324 57134
rect 109084 56866 109324 56898
rect 118084 57454 118324 57486
rect 118084 57218 118086 57454
rect 118322 57218 118324 57454
rect 118084 57134 118324 57218
rect 118084 56898 118086 57134
rect 118322 56898 118324 57134
rect 118084 56866 118324 56898
rect 127084 57454 127324 57486
rect 127084 57218 127086 57454
rect 127322 57218 127324 57454
rect 127084 57134 127324 57218
rect 127084 56898 127086 57134
rect 127322 56898 127324 57134
rect 127084 56866 127324 56898
rect 136084 57454 136324 57486
rect 136084 57218 136086 57454
rect 136322 57218 136324 57454
rect 136084 57134 136324 57218
rect 136084 56898 136086 57134
rect 136322 56898 136324 57134
rect 136084 56866 136324 56898
rect 145084 57454 145324 57486
rect 145084 57218 145086 57454
rect 145322 57218 145324 57454
rect 145084 57134 145324 57218
rect 145084 56898 145086 57134
rect 145322 56898 145324 57134
rect 145084 56866 145324 56898
rect 147646 57454 147886 57486
rect 147646 57218 147648 57454
rect 147884 57218 147886 57454
rect 147646 57134 147886 57218
rect 147646 56898 147648 57134
rect 147884 56898 147886 57134
rect 147646 56866 147886 56898
rect 149298 57454 149538 57486
rect 149298 57218 149300 57454
rect 149536 57218 149538 57454
rect 149298 57134 149538 57218
rect 149298 56898 149300 57134
rect 149536 56898 149538 57134
rect 149298 56866 149538 56898
rect 150104 57454 150344 57486
rect 150104 57218 150106 57454
rect 150342 57218 150344 57454
rect 150104 57134 150344 57218
rect 150104 56898 150106 57134
rect 150342 56898 150344 57134
rect 150104 56866 150344 56898
rect 159104 57454 159344 57486
rect 159104 57218 159106 57454
rect 159342 57218 159344 57454
rect 159104 57134 159344 57218
rect 159104 56898 159106 57134
rect 159342 56898 159344 57134
rect 159104 56866 159344 56898
rect 168104 57454 168344 57486
rect 168104 57218 168106 57454
rect 168342 57218 168344 57454
rect 168104 57134 168344 57218
rect 168104 56898 168106 57134
rect 168342 56898 168344 57134
rect 168104 56866 168344 56898
rect 177104 57454 177344 57486
rect 177104 57218 177106 57454
rect 177342 57218 177344 57454
rect 177104 57134 177344 57218
rect 177104 56898 177106 57134
rect 177342 56898 177344 57134
rect 177104 56866 177344 56898
rect 186104 57454 186344 57486
rect 186104 57218 186106 57454
rect 186342 57218 186344 57454
rect 186104 57134 186344 57218
rect 186104 56898 186106 57134
rect 186342 56898 186344 57134
rect 186104 56866 186344 56898
rect 188666 57454 188906 57486
rect 188666 57218 188668 57454
rect 188904 57218 188906 57454
rect 188666 57134 188906 57218
rect 188666 56898 188668 57134
rect 188904 56898 188906 57134
rect 188666 56866 188906 56898
rect 190318 57454 190558 57486
rect 190318 57218 190320 57454
rect 190556 57218 190558 57454
rect 190318 57134 190558 57218
rect 190318 56898 190320 57134
rect 190556 56898 190558 57134
rect 190318 56866 190558 56898
rect 191124 57454 191364 57486
rect 191124 57218 191126 57454
rect 191362 57218 191364 57454
rect 191124 57134 191364 57218
rect 191124 56898 191126 57134
rect 191362 56898 191364 57134
rect 191124 56866 191364 56898
rect 200124 57454 200364 57486
rect 200124 57218 200126 57454
rect 200362 57218 200364 57454
rect 200124 57134 200364 57218
rect 200124 56898 200126 57134
rect 200362 56898 200364 57134
rect 200124 56866 200364 56898
rect 209124 57454 209364 57486
rect 209124 57218 209126 57454
rect 209362 57218 209364 57454
rect 209124 57134 209364 57218
rect 209124 56898 209126 57134
rect 209362 56898 209364 57134
rect 209124 56866 209364 56898
rect 218124 57454 218364 57486
rect 218124 57218 218126 57454
rect 218362 57218 218364 57454
rect 218124 57134 218364 57218
rect 218124 56898 218126 57134
rect 218362 56898 218364 57134
rect 218124 56866 218364 56898
rect 227124 57454 227364 57486
rect 227124 57218 227126 57454
rect 227362 57218 227364 57454
rect 227124 57134 227364 57218
rect 227124 56898 227126 57134
rect 227362 56898 227364 57134
rect 227124 56866 227364 56898
rect 229686 57454 229926 57486
rect 229686 57218 229688 57454
rect 229924 57218 229926 57454
rect 229686 57134 229926 57218
rect 229686 56898 229688 57134
rect 229924 56898 229926 57134
rect 229686 56866 229926 56898
rect 230338 57454 230578 57486
rect 230338 57218 230340 57454
rect 230576 57218 230578 57454
rect 230338 57134 230578 57218
rect 230338 56898 230340 57134
rect 230576 56898 230578 57134
rect 230338 56866 230578 56898
rect 231144 57454 231384 57486
rect 231144 57218 231146 57454
rect 231382 57218 231384 57454
rect 231144 57134 231384 57218
rect 231144 56898 231146 57134
rect 231382 56898 231384 57134
rect 231144 56866 231384 56898
rect 240144 57454 240384 57486
rect 240144 57218 240146 57454
rect 240382 57218 240384 57454
rect 240144 57134 240384 57218
rect 240144 56898 240146 57134
rect 240382 56898 240384 57134
rect 240144 56866 240384 56898
rect 249144 57454 249384 57486
rect 249144 57218 249146 57454
rect 249382 57218 249384 57454
rect 249144 57134 249384 57218
rect 249144 56898 249146 57134
rect 249382 56898 249384 57134
rect 249144 56866 249384 56898
rect 258144 57454 258384 57486
rect 258144 57218 258146 57454
rect 258382 57218 258384 57454
rect 258144 57134 258384 57218
rect 258144 56898 258146 57134
rect 258382 56898 258384 57134
rect 258144 56866 258384 56898
rect 267144 57454 267384 57486
rect 267144 57218 267146 57454
rect 267382 57218 267384 57454
rect 267144 57134 267384 57218
rect 267144 56898 267146 57134
rect 267382 56898 267384 57134
rect 267144 56866 267384 56898
rect 269706 57454 269946 57486
rect 269706 57218 269708 57454
rect 269944 57218 269946 57454
rect 269706 57134 269946 57218
rect 269706 56898 269708 57134
rect 269944 56898 269946 57134
rect 269706 56866 269946 56898
rect 270358 57454 270598 57486
rect 270358 57218 270360 57454
rect 270596 57218 270598 57454
rect 270358 57134 270598 57218
rect 270358 56898 270360 57134
rect 270596 56898 270598 57134
rect 270358 56866 270598 56898
rect 271164 57454 271404 57486
rect 271164 57218 271166 57454
rect 271402 57218 271404 57454
rect 271164 57134 271404 57218
rect 271164 56898 271166 57134
rect 271402 56898 271404 57134
rect 271164 56866 271404 56898
rect 280164 57454 280404 57486
rect 280164 57218 280166 57454
rect 280402 57218 280404 57454
rect 280164 57134 280404 57218
rect 280164 56898 280166 57134
rect 280402 56898 280404 57134
rect 280164 56866 280404 56898
rect 289164 57454 289404 57486
rect 289164 57218 289166 57454
rect 289402 57218 289404 57454
rect 289164 57134 289404 57218
rect 289164 56898 289166 57134
rect 289402 56898 289404 57134
rect 289164 56866 289404 56898
rect 298164 57454 298404 57486
rect 298164 57218 298166 57454
rect 298402 57218 298404 57454
rect 298164 57134 298404 57218
rect 298164 56898 298166 57134
rect 298402 56898 298404 57134
rect 298164 56866 298404 56898
rect 307164 57454 307404 57486
rect 307164 57218 307166 57454
rect 307402 57218 307404 57454
rect 307164 57134 307404 57218
rect 307164 56898 307166 57134
rect 307402 56898 307404 57134
rect 307164 56866 307404 56898
rect 309726 57454 309966 57486
rect 309726 57218 309728 57454
rect 309964 57218 309966 57454
rect 309726 57134 309966 57218
rect 309726 56898 309728 57134
rect 309964 56898 309966 57134
rect 309726 56866 309966 56898
rect 311378 57454 311618 57486
rect 311378 57218 311380 57454
rect 311616 57218 311618 57454
rect 311378 57134 311618 57218
rect 311378 56898 311380 57134
rect 311616 56898 311618 57134
rect 311378 56866 311618 56898
rect 312184 57454 312424 57486
rect 312184 57218 312186 57454
rect 312422 57218 312424 57454
rect 312184 57134 312424 57218
rect 312184 56898 312186 57134
rect 312422 56898 312424 57134
rect 312184 56866 312424 56898
rect 321184 57454 321424 57486
rect 321184 57218 321186 57454
rect 321422 57218 321424 57454
rect 321184 57134 321424 57218
rect 321184 56898 321186 57134
rect 321422 56898 321424 57134
rect 321184 56866 321424 56898
rect 330184 57454 330424 57486
rect 330184 57218 330186 57454
rect 330422 57218 330424 57454
rect 330184 57134 330424 57218
rect 330184 56898 330186 57134
rect 330422 56898 330424 57134
rect 330184 56866 330424 56898
rect 339184 57454 339424 57486
rect 339184 57218 339186 57454
rect 339422 57218 339424 57454
rect 339184 57134 339424 57218
rect 339184 56898 339186 57134
rect 339422 56898 339424 57134
rect 339184 56866 339424 56898
rect 348184 57454 348424 57486
rect 348184 57218 348186 57454
rect 348422 57218 348424 57454
rect 348184 57134 348424 57218
rect 348184 56898 348186 57134
rect 348422 56898 348424 57134
rect 348184 56866 348424 56898
rect 350746 57454 350986 57486
rect 350746 57218 350748 57454
rect 350984 57218 350986 57454
rect 350746 57134 350986 57218
rect 350746 56898 350748 57134
rect 350984 56898 350986 57134
rect 350746 56866 350986 56898
rect 352398 57454 352638 57486
rect 352398 57218 352400 57454
rect 352636 57218 352638 57454
rect 352398 57134 352638 57218
rect 352398 56898 352400 57134
rect 352636 56898 352638 57134
rect 352398 56866 352638 56898
rect 353204 57454 353444 57486
rect 353204 57218 353206 57454
rect 353442 57218 353444 57454
rect 353204 57134 353444 57218
rect 353204 56898 353206 57134
rect 353442 56898 353444 57134
rect 353204 56866 353444 56898
rect 362204 57454 362444 57486
rect 362204 57218 362206 57454
rect 362442 57218 362444 57454
rect 362204 57134 362444 57218
rect 362204 56898 362206 57134
rect 362442 56898 362444 57134
rect 362204 56866 362444 56898
rect 371204 57454 371444 57486
rect 371204 57218 371206 57454
rect 371442 57218 371444 57454
rect 371204 57134 371444 57218
rect 371204 56898 371206 57134
rect 371442 56898 371444 57134
rect 371204 56866 371444 56898
rect 380204 57454 380444 57486
rect 380204 57218 380206 57454
rect 380442 57218 380444 57454
rect 380204 57134 380444 57218
rect 380204 56898 380206 57134
rect 380442 56898 380444 57134
rect 380204 56866 380444 56898
rect 389204 57454 389444 57486
rect 389204 57218 389206 57454
rect 389442 57218 389444 57454
rect 389204 57134 389444 57218
rect 389204 56898 389206 57134
rect 389442 56898 389444 57134
rect 389204 56866 389444 56898
rect 391766 57454 392006 57486
rect 391766 57218 391768 57454
rect 392004 57218 392006 57454
rect 391766 57134 392006 57218
rect 391766 56898 391768 57134
rect 392004 56898 392006 57134
rect 391766 56866 392006 56898
rect 392418 57454 392658 57486
rect 392418 57218 392420 57454
rect 392656 57218 392658 57454
rect 392418 57134 392658 57218
rect 392418 56898 392420 57134
rect 392656 56898 392658 57134
rect 392418 56866 392658 56898
rect 393224 57454 393464 57486
rect 393224 57218 393226 57454
rect 393462 57218 393464 57454
rect 393224 57134 393464 57218
rect 393224 56898 393226 57134
rect 393462 56898 393464 57134
rect 393224 56866 393464 56898
rect 402224 57454 402464 57486
rect 402224 57218 402226 57454
rect 402462 57218 402464 57454
rect 402224 57134 402464 57218
rect 402224 56898 402226 57134
rect 402462 56898 402464 57134
rect 402224 56866 402464 56898
rect 411224 57454 411464 57486
rect 411224 57218 411226 57454
rect 411462 57218 411464 57454
rect 411224 57134 411464 57218
rect 411224 56898 411226 57134
rect 411462 56898 411464 57134
rect 411224 56866 411464 56898
rect 420224 57454 420464 57486
rect 420224 57218 420226 57454
rect 420462 57218 420464 57454
rect 420224 57134 420464 57218
rect 420224 56898 420226 57134
rect 420462 56898 420464 57134
rect 420224 56866 420464 56898
rect 429224 57454 429464 57486
rect 429224 57218 429226 57454
rect 429462 57218 429464 57454
rect 429224 57134 429464 57218
rect 429224 56898 429226 57134
rect 429462 56898 429464 57134
rect 429224 56866 429464 56898
rect 431786 57454 432026 57486
rect 431786 57218 431788 57454
rect 432024 57218 432026 57454
rect 431786 57134 432026 57218
rect 431786 56898 431788 57134
rect 432024 56898 432026 57134
rect 431786 56866 432026 56898
rect 432438 57454 432678 57486
rect 432438 57218 432440 57454
rect 432676 57218 432678 57454
rect 432438 57134 432678 57218
rect 432438 56898 432440 57134
rect 432676 56898 432678 57134
rect 432438 56866 432678 56898
rect 433244 57454 433484 57486
rect 433244 57218 433246 57454
rect 433482 57218 433484 57454
rect 433244 57134 433484 57218
rect 433244 56898 433246 57134
rect 433482 56898 433484 57134
rect 433244 56866 433484 56898
rect 442244 57454 442484 57486
rect 442244 57218 442246 57454
rect 442482 57218 442484 57454
rect 442244 57134 442484 57218
rect 442244 56898 442246 57134
rect 442482 56898 442484 57134
rect 442244 56866 442484 56898
rect 451244 57454 451484 57486
rect 451244 57218 451246 57454
rect 451482 57218 451484 57454
rect 451244 57134 451484 57218
rect 451244 56898 451246 57134
rect 451482 56898 451484 57134
rect 451244 56866 451484 56898
rect 460244 57454 460484 57486
rect 460244 57218 460246 57454
rect 460482 57218 460484 57454
rect 460244 57134 460484 57218
rect 460244 56898 460246 57134
rect 460482 56898 460484 57134
rect 460244 56866 460484 56898
rect 469244 57454 469484 57486
rect 469244 57218 469246 57454
rect 469482 57218 469484 57454
rect 469244 57134 469484 57218
rect 469244 56898 469246 57134
rect 469482 56898 469484 57134
rect 469244 56866 469484 56898
rect 471806 57454 472046 57486
rect 471806 57218 471808 57454
rect 472044 57218 472046 57454
rect 471806 57134 472046 57218
rect 471806 56898 471808 57134
rect 472044 56898 472046 57134
rect 471806 56866 472046 56898
rect 472458 57454 472698 57486
rect 472458 57218 472460 57454
rect 472696 57218 472698 57454
rect 472458 57134 472698 57218
rect 472458 56898 472460 57134
rect 472696 56898 472698 57134
rect 472458 56866 472698 56898
rect 473264 57454 473504 57486
rect 473264 57218 473266 57454
rect 473502 57218 473504 57454
rect 473264 57134 473504 57218
rect 473264 56898 473266 57134
rect 473502 56898 473504 57134
rect 473264 56866 473504 56898
rect 482264 57454 482504 57486
rect 482264 57218 482266 57454
rect 482502 57218 482504 57454
rect 482264 57134 482504 57218
rect 482264 56898 482266 57134
rect 482502 56898 482504 57134
rect 482264 56866 482504 56898
rect 491264 57454 491504 57486
rect 491264 57218 491266 57454
rect 491502 57218 491504 57454
rect 491264 57134 491504 57218
rect 491264 56898 491266 57134
rect 491502 56898 491504 57134
rect 491264 56866 491504 56898
rect 500264 57454 500504 57486
rect 500264 57218 500266 57454
rect 500502 57218 500504 57454
rect 500264 57134 500504 57218
rect 500264 56898 500266 57134
rect 500502 56898 500504 57134
rect 500264 56866 500504 56898
rect 509264 57454 509504 57486
rect 509264 57218 509266 57454
rect 509502 57218 509504 57454
rect 509264 57134 509504 57218
rect 509264 56898 509266 57134
rect 509502 56898 509504 57134
rect 509264 56866 509504 56898
rect 511826 57454 512066 57486
rect 511826 57218 511828 57454
rect 512064 57218 512066 57454
rect 511826 57134 512066 57218
rect 511826 56898 511828 57134
rect 512064 56898 512066 57134
rect 511826 56866 512066 56898
rect 512478 57454 512718 57486
rect 512478 57218 512480 57454
rect 512716 57218 512718 57454
rect 512478 57134 512718 57218
rect 512478 56898 512480 57134
rect 512716 56898 512718 57134
rect 512478 56866 512718 56898
rect 513284 57454 513524 57486
rect 513284 57218 513286 57454
rect 513522 57218 513524 57454
rect 513284 57134 513524 57218
rect 513284 56898 513286 57134
rect 513522 56898 513524 57134
rect 513284 56866 513524 56898
rect 522284 57454 522524 57486
rect 522284 57218 522286 57454
rect 522522 57218 522524 57454
rect 522284 57134 522524 57218
rect 522284 56898 522286 57134
rect 522522 56898 522524 57134
rect 522284 56866 522524 56898
rect 531284 57454 531524 57486
rect 531284 57218 531286 57454
rect 531522 57218 531524 57454
rect 531284 57134 531524 57218
rect 531284 56898 531286 57134
rect 531522 56898 531524 57134
rect 531284 56866 531524 56898
rect 540284 57454 540524 57486
rect 540284 57218 540286 57454
rect 540522 57218 540524 57454
rect 540284 57134 540524 57218
rect 540284 56898 540286 57134
rect 540522 56898 540524 57134
rect 540284 56866 540524 56898
rect 549284 57454 549524 57486
rect 549284 57218 549286 57454
rect 549522 57218 549524 57454
rect 549284 57134 549524 57218
rect 549284 56898 549286 57134
rect 549522 56898 549524 57134
rect 549284 56866 549524 56898
rect 551846 57454 552086 57486
rect 551846 57218 551848 57454
rect 552084 57218 552086 57454
rect 551846 57134 552086 57218
rect 551846 56898 551848 57134
rect 552084 56898 552086 57134
rect 551846 56866 552086 56898
rect 552498 57454 552738 57486
rect 552498 57218 552500 57454
rect 552736 57218 552738 57454
rect 552498 57134 552738 57218
rect 552498 56898 552500 57134
rect 552736 56898 552738 57134
rect 552498 56866 552738 56898
rect 553304 57454 553544 57486
rect 553304 57218 553306 57454
rect 553542 57218 553544 57454
rect 553304 57134 553544 57218
rect 553304 56898 553306 57134
rect 553542 56898 553544 57134
rect 553304 56866 553544 56898
rect 562304 57454 562544 57486
rect 562304 57218 562306 57454
rect 562542 57218 562544 57454
rect 562304 57134 562544 57218
rect 562304 56898 562306 57134
rect 562542 56898 562544 57134
rect 562304 56866 562544 56898
rect 571304 57454 571544 57486
rect 571304 57218 571306 57454
rect 571542 57218 571544 57454
rect 571304 57134 571544 57218
rect 571304 56898 571306 57134
rect 571542 56898 571544 57134
rect 571304 56866 571544 56898
rect 573834 57454 574074 57486
rect 573834 57218 573836 57454
rect 574072 57218 574074 57454
rect 573834 57134 574074 57218
rect 573834 56898 573836 57134
rect 574072 56898 574074 57134
rect 573834 56866 574074 56898
rect 579288 57454 579888 57486
rect 579288 57218 579470 57454
rect 579706 57218 579888 57454
rect 579288 57134 579888 57218
rect 579288 56898 579470 57134
rect 579706 56898 579888 57134
rect 579288 56866 579888 56898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect 5200 39454 5800 39486
rect 5200 39218 5382 39454
rect 5618 39218 5800 39454
rect 5200 39134 5800 39218
rect 5200 38898 5382 39134
rect 5618 38898 5800 39134
rect 5200 38866 5800 38898
rect 578488 39454 579088 39486
rect 578488 39218 578670 39454
rect 578906 39218 579088 39454
rect 578488 39134 579088 39218
rect 578488 38898 578670 39134
rect 578906 38898 579088 39134
rect 578488 38866 579088 38898
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 3454 2414 28000
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 7174 6134 28000
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 10894 9854 28000
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 14614 13574 28000
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 21454 20414 28000
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 25174 24134 28000
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 -5146 27854 28000
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 28000
rect 37794 3454 38414 28000
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 7174 42134 28000
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 10894 45854 28000
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 14614 49574 28000
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 21454 56414 28000
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 28000
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 -5146 63854 28000
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 28000
rect 73794 3454 74414 28000
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 7174 78134 28000
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 10894 81854 28000
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 14614 85574 28000
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 21454 92414 28000
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 28000
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 -5146 99854 28000
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 28000
rect 109794 3454 110414 28000
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 7174 114134 28000
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 10894 117854 28000
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 14614 121574 28000
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 21454 128414 28000
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 28000
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 -5146 135854 28000
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 28000
rect 145794 3454 146414 28000
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 7174 150134 28000
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 10894 153854 28000
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 14614 157574 28000
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 21454 164414 28000
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 28000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 -5146 171854 28000
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 28000
rect 181794 3454 182414 28000
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 7174 186134 28000
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 10894 189854 28000
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 14614 193574 28000
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 21454 200414 28000
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 28000
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 -5146 207854 28000
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 28000
rect 217794 3454 218414 28000
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 7174 222134 28000
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 10894 225854 28000
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 14614 229574 28000
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 21454 236414 28000
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 28000
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 -5146 243854 28000
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 28000
rect 253794 3454 254414 28000
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 7174 258134 28000
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 10894 261854 28000
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 14614 265574 28000
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 28000
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 28000
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 -5146 279854 28000
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 28000
rect 289794 3454 290414 28000
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 7174 294134 28000
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 10894 297854 28000
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 14614 301574 28000
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 21454 308414 28000
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 28000
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 -5146 315854 28000
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 28000
rect 325794 3454 326414 28000
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 7174 330134 28000
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 10894 333854 28000
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 14614 337574 28000
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 21454 344414 28000
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 28000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 -5146 351854 28000
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 28000
rect 361794 3454 362414 28000
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 7174 366134 28000
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 10894 369854 28000
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 14614 373574 28000
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 21454 380414 28000
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 28000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 -5146 387854 28000
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 28000
rect 397794 3454 398414 28000
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 7174 402134 28000
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 10894 405854 28000
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 14614 409574 28000
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 21454 416414 28000
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 28000
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 -5146 423854 28000
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 28000
rect 433794 3454 434414 28000
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 7174 438134 28000
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 10894 441854 28000
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 14614 445574 28000
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 21454 452414 28000
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 28000
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 -5146 459854 28000
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 28000
rect 469794 3454 470414 28000
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 7174 474134 28000
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 10894 477854 28000
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 14614 481574 28000
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 21454 488414 28000
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 25174 492134 28000
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 -5146 495854 28000
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 28000
rect 505794 3454 506414 28000
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 7174 510134 28000
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 10894 513854 28000
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 14614 517574 28000
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 21454 524414 28000
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 25174 528134 28000
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 -5146 531854 28000
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 28000
rect 541794 3454 542414 28000
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 7174 546134 28000
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 10894 549854 28000
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 14614 553574 28000
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 21454 560414 28000
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 25174 564134 28000
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 -5146 567854 28000
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 28000
rect 577794 3454 578414 28000
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 7174 582134 28000
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 4582 669218 4818 669454
rect 4582 668898 4818 669134
rect 127058 669218 127294 669454
rect 127058 668898 127294 669134
rect 140296 669218 140532 669454
rect 140296 668898 140532 669134
rect 147648 669218 147884 669454
rect 147648 668898 147884 669134
rect 190320 669218 190556 669454
rect 190320 668898 190556 669134
rect 229688 669218 229924 669454
rect 229688 668898 229924 669134
rect 432440 669218 432676 669454
rect 432440 668898 432676 669134
rect 439792 669218 440028 669454
rect 439792 668898 440028 669134
rect 457010 669218 457246 669454
rect 457010 668898 457246 669134
rect 579470 669218 579706 669454
rect 579470 668898 579706 669134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect 5382 651218 5618 651454
rect 5382 650898 5618 651134
rect 127458 651218 127694 651454
rect 127458 650898 127694 651134
rect 140656 651218 140892 651454
rect 140656 650898 140892 651134
rect 147288 651218 147524 651454
rect 147288 650898 147524 651134
rect 149660 651218 149896 651454
rect 149660 650898 149896 651134
rect 188308 651218 188544 651454
rect 188308 650898 188544 651134
rect 190680 651218 190916 651454
rect 190680 650898 190916 651134
rect 229328 651218 229564 651454
rect 229328 650898 229564 651134
rect 230700 651218 230936 651454
rect 230700 650898 230936 651134
rect 269348 651218 269584 651454
rect 269348 650898 269584 651134
rect 270720 651218 270956 651454
rect 270720 650898 270956 651134
rect 309368 651218 309604 651454
rect 309368 650898 309604 651134
rect 310564 651218 310800 651454
rect 310564 650898 310800 651134
rect 311740 651218 311976 651454
rect 311740 650898 311976 651134
rect 350388 651218 350624 651454
rect 350388 650898 350624 651134
rect 352760 651218 352996 651454
rect 352760 650898 352996 651134
rect 391408 651218 391644 651454
rect 391408 650898 391644 651134
rect 392780 651218 393016 651454
rect 392780 650898 393016 651134
rect 431428 651218 431664 651454
rect 431428 650898 431664 651134
rect 432800 651218 433036 651454
rect 432800 650898 433036 651134
rect 439432 651218 439668 651454
rect 439432 650898 439668 651134
rect 456610 651218 456846 651454
rect 456610 650898 456846 651134
rect 578670 651218 578906 651454
rect 578670 650898 578906 651134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 4582 633218 4818 633454
rect 4582 632898 4818 633134
rect 12352 633218 12588 633454
rect 12352 632898 12588 633134
rect 107416 633218 107652 633454
rect 107416 632898 107652 633134
rect 127058 633218 127294 633454
rect 127058 632898 127294 633134
rect 140296 633218 140532 633454
rect 140296 632898 140532 633134
rect 141102 633218 141338 633454
rect 141102 632898 141338 633134
rect 147648 633218 147884 633454
rect 147648 632898 147884 633134
rect 149300 633218 149536 633454
rect 149300 632898 149536 633134
rect 150106 633218 150342 633454
rect 150106 632898 150342 633134
rect 159106 633218 159342 633454
rect 159106 632898 159342 633134
rect 168106 633218 168342 633454
rect 168106 632898 168342 633134
rect 177106 633218 177342 633454
rect 177106 632898 177342 633134
rect 186106 633218 186342 633454
rect 186106 632898 186342 633134
rect 188668 633218 188904 633454
rect 188668 632898 188904 633134
rect 190320 633218 190556 633454
rect 190320 632898 190556 633134
rect 191126 633218 191362 633454
rect 191126 632898 191362 633134
rect 200126 633218 200362 633454
rect 200126 632898 200362 633134
rect 209126 633218 209362 633454
rect 209126 632898 209362 633134
rect 218126 633218 218362 633454
rect 218126 632898 218362 633134
rect 227126 633218 227362 633454
rect 227126 632898 227362 633134
rect 229688 633218 229924 633454
rect 229688 632898 229924 633134
rect 230340 633218 230576 633454
rect 230340 632898 230576 633134
rect 231146 633218 231382 633454
rect 231146 632898 231382 633134
rect 240146 633218 240382 633454
rect 240146 632898 240382 633134
rect 249146 633218 249382 633454
rect 249146 632898 249382 633134
rect 258146 633218 258382 633454
rect 258146 632898 258382 633134
rect 267146 633218 267382 633454
rect 267146 632898 267382 633134
rect 269708 633218 269944 633454
rect 269708 632898 269944 633134
rect 270360 633218 270596 633454
rect 270360 632898 270596 633134
rect 271166 633218 271402 633454
rect 271166 632898 271402 633134
rect 280166 633218 280402 633454
rect 280166 632898 280402 633134
rect 289166 633218 289402 633454
rect 289166 632898 289402 633134
rect 298166 633218 298402 633454
rect 298166 632898 298402 633134
rect 307166 633218 307402 633454
rect 307166 632898 307402 633134
rect 309728 633218 309964 633454
rect 309728 632898 309964 633134
rect 311380 633218 311616 633454
rect 311380 632898 311616 633134
rect 312186 633218 312422 633454
rect 312186 632898 312422 633134
rect 321186 633218 321422 633454
rect 321186 632898 321422 633134
rect 330186 633218 330422 633454
rect 330186 632898 330422 633134
rect 339186 633218 339422 633454
rect 339186 632898 339422 633134
rect 348186 633218 348422 633454
rect 348186 632898 348422 633134
rect 350748 633218 350984 633454
rect 350748 632898 350984 633134
rect 352400 633218 352636 633454
rect 352400 632898 352636 633134
rect 353206 633218 353442 633454
rect 353206 632898 353442 633134
rect 362206 633218 362442 633454
rect 362206 632898 362442 633134
rect 371206 633218 371442 633454
rect 371206 632898 371442 633134
rect 380206 633218 380442 633454
rect 380206 632898 380442 633134
rect 389206 633218 389442 633454
rect 389206 632898 389442 633134
rect 391768 633218 392004 633454
rect 391768 632898 392004 633134
rect 392420 633218 392656 633454
rect 392420 632898 392656 633134
rect 393226 633218 393462 633454
rect 393226 632898 393462 633134
rect 402226 633218 402462 633454
rect 402226 632898 402462 633134
rect 411226 633218 411462 633454
rect 411226 632898 411462 633134
rect 420226 633218 420462 633454
rect 420226 632898 420462 633134
rect 429226 633218 429462 633454
rect 429226 632898 429462 633134
rect 431788 633218 432024 633454
rect 431788 632898 432024 633134
rect 432440 633218 432676 633454
rect 432440 632898 432676 633134
rect 433246 633218 433482 633454
rect 433246 632898 433482 633134
rect 439792 633218 440028 633454
rect 439792 632898 440028 633134
rect 457010 633218 457246 633454
rect 457010 632898 457246 633134
rect 476652 633218 476888 633454
rect 476652 632898 476888 633134
rect 571716 633218 571952 633454
rect 571716 632898 571952 633134
rect 579470 633218 579706 633454
rect 579470 632898 579706 633134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect 5382 615218 5618 615454
rect 5382 614898 5618 615134
rect 13032 615218 13268 615454
rect 13032 614898 13268 615134
rect 106736 615218 106972 615454
rect 106736 614898 106972 615134
rect 127458 615218 127694 615454
rect 127458 614898 127694 615134
rect 140656 615218 140892 615454
rect 140656 614898 140892 615134
rect 141502 615218 141738 615454
rect 141502 614898 141738 615134
rect 147288 615218 147524 615454
rect 147288 614898 147524 615134
rect 149660 615218 149896 615454
rect 149660 614898 149896 615134
rect 150506 615218 150742 615454
rect 150506 614898 150742 615134
rect 159506 615218 159742 615454
rect 159506 614898 159742 615134
rect 168506 615218 168742 615454
rect 168506 614898 168742 615134
rect 177506 615218 177742 615454
rect 177506 614898 177742 615134
rect 186506 615218 186742 615454
rect 186506 614898 186742 615134
rect 188308 615218 188544 615454
rect 188308 614898 188544 615134
rect 190680 615218 190916 615454
rect 190680 614898 190916 615134
rect 191526 615218 191762 615454
rect 191526 614898 191762 615134
rect 200526 615218 200762 615454
rect 200526 614898 200762 615134
rect 209526 615218 209762 615454
rect 209526 614898 209762 615134
rect 218526 615218 218762 615454
rect 218526 614898 218762 615134
rect 227526 615218 227762 615454
rect 227526 614898 227762 615134
rect 229328 615218 229564 615454
rect 229328 614898 229564 615134
rect 230700 615218 230936 615454
rect 230700 614898 230936 615134
rect 231546 615218 231782 615454
rect 231546 614898 231782 615134
rect 240546 615218 240782 615454
rect 240546 614898 240782 615134
rect 249546 615218 249782 615454
rect 249546 614898 249782 615134
rect 258546 615218 258782 615454
rect 258546 614898 258782 615134
rect 267546 615218 267782 615454
rect 267546 614898 267782 615134
rect 269348 615218 269584 615454
rect 269348 614898 269584 615134
rect 270720 615218 270956 615454
rect 270720 614898 270956 615134
rect 271566 615218 271802 615454
rect 271566 614898 271802 615134
rect 280566 615218 280802 615454
rect 280566 614898 280802 615134
rect 289566 615218 289802 615454
rect 289566 614898 289802 615134
rect 298566 615218 298802 615454
rect 298566 614898 298802 615134
rect 307566 615218 307802 615454
rect 307566 614898 307802 615134
rect 309368 615218 309604 615454
rect 309368 614898 309604 615134
rect 311740 615218 311976 615454
rect 311740 614898 311976 615134
rect 312586 615218 312822 615454
rect 312586 614898 312822 615134
rect 321586 615218 321822 615454
rect 321586 614898 321822 615134
rect 330586 615218 330822 615454
rect 330586 614898 330822 615134
rect 339586 615218 339822 615454
rect 339586 614898 339822 615134
rect 348586 615218 348822 615454
rect 348586 614898 348822 615134
rect 350388 615218 350624 615454
rect 350388 614898 350624 615134
rect 352760 615218 352996 615454
rect 352760 614898 352996 615134
rect 353606 615218 353842 615454
rect 353606 614898 353842 615134
rect 362606 615218 362842 615454
rect 362606 614898 362842 615134
rect 371606 615218 371842 615454
rect 371606 614898 371842 615134
rect 380606 615218 380842 615454
rect 380606 614898 380842 615134
rect 389606 615218 389842 615454
rect 389606 614898 389842 615134
rect 391408 615218 391644 615454
rect 391408 614898 391644 615134
rect 392780 615218 393016 615454
rect 392780 614898 393016 615134
rect 393626 615218 393862 615454
rect 393626 614898 393862 615134
rect 402626 615218 402862 615454
rect 402626 614898 402862 615134
rect 411626 615218 411862 615454
rect 411626 614898 411862 615134
rect 420626 615218 420862 615454
rect 420626 614898 420862 615134
rect 429626 615218 429862 615454
rect 429626 614898 429862 615134
rect 431428 615218 431664 615454
rect 431428 614898 431664 615134
rect 432800 615218 433036 615454
rect 432800 614898 433036 615134
rect 433646 615218 433882 615454
rect 433646 614898 433882 615134
rect 439432 615218 439668 615454
rect 439432 614898 439668 615134
rect 456610 615218 456846 615454
rect 456610 614898 456846 615134
rect 477332 615218 477568 615454
rect 477332 614898 477568 615134
rect 571036 615218 571272 615454
rect 571036 614898 571272 615134
rect 578670 615218 578906 615454
rect 578670 614898 578906 615134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 4582 597218 4818 597454
rect 4582 596898 4818 597134
rect 12352 597218 12588 597454
rect 12352 596898 12588 597134
rect 107416 597218 107652 597454
rect 107416 596898 107652 597134
rect 127058 597218 127294 597454
rect 127058 596898 127294 597134
rect 140296 597218 140532 597454
rect 140296 596898 140532 597134
rect 141102 597218 141338 597454
rect 141102 596898 141338 597134
rect 147648 597218 147884 597454
rect 147648 596898 147884 597134
rect 149300 597218 149536 597454
rect 149300 596898 149536 597134
rect 150106 597218 150342 597454
rect 150106 596898 150342 597134
rect 159106 597218 159342 597454
rect 159106 596898 159342 597134
rect 168106 597218 168342 597454
rect 168106 596898 168342 597134
rect 177106 597218 177342 597454
rect 177106 596898 177342 597134
rect 186106 597218 186342 597454
rect 186106 596898 186342 597134
rect 188668 597218 188904 597454
rect 188668 596898 188904 597134
rect 189768 597218 190004 597454
rect 189768 596898 190004 597134
rect 190320 597218 190556 597454
rect 190320 596898 190556 597134
rect 191126 597218 191362 597454
rect 191126 596898 191362 597134
rect 200126 597218 200362 597454
rect 200126 596898 200362 597134
rect 209126 597218 209362 597454
rect 209126 596898 209362 597134
rect 218126 597218 218362 597454
rect 218126 596898 218362 597134
rect 227126 597218 227362 597454
rect 227126 596898 227362 597134
rect 229688 597218 229924 597454
rect 229688 596898 229924 597134
rect 230340 597218 230576 597454
rect 230340 596898 230576 597134
rect 231146 597218 231382 597454
rect 231146 596898 231382 597134
rect 240146 597218 240382 597454
rect 240146 596898 240382 597134
rect 249146 597218 249382 597454
rect 249146 596898 249382 597134
rect 258146 597218 258382 597454
rect 258146 596898 258382 597134
rect 267146 597218 267382 597454
rect 267146 596898 267382 597134
rect 269708 597218 269944 597454
rect 269708 596898 269944 597134
rect 270360 597218 270596 597454
rect 270360 596898 270596 597134
rect 271166 597218 271402 597454
rect 271166 596898 271402 597134
rect 280166 597218 280402 597454
rect 280166 596898 280402 597134
rect 289166 597218 289402 597454
rect 289166 596898 289402 597134
rect 298166 597218 298402 597454
rect 298166 596898 298402 597134
rect 307166 597218 307402 597454
rect 307166 596898 307402 597134
rect 309728 597218 309964 597454
rect 309728 596898 309964 597134
rect 311380 597218 311616 597454
rect 311380 596898 311616 597134
rect 312186 597218 312422 597454
rect 312186 596898 312422 597134
rect 321186 597218 321422 597454
rect 321186 596898 321422 597134
rect 330186 597218 330422 597454
rect 330186 596898 330422 597134
rect 339186 597218 339422 597454
rect 339186 596898 339422 597134
rect 348186 597218 348422 597454
rect 348186 596898 348422 597134
rect 350748 597218 350984 597454
rect 350748 596898 350984 597134
rect 352400 597218 352636 597454
rect 352400 596898 352636 597134
rect 353206 597218 353442 597454
rect 353206 596898 353442 597134
rect 362206 597218 362442 597454
rect 362206 596898 362442 597134
rect 371206 597218 371442 597454
rect 371206 596898 371442 597134
rect 380206 597218 380442 597454
rect 380206 596898 380442 597134
rect 389206 597218 389442 597454
rect 389206 596898 389442 597134
rect 391768 597218 392004 597454
rect 391768 596898 392004 597134
rect 392420 597218 392656 597454
rect 392420 596898 392656 597134
rect 393226 597218 393462 597454
rect 393226 596898 393462 597134
rect 402226 597218 402462 597454
rect 402226 596898 402462 597134
rect 411226 597218 411462 597454
rect 411226 596898 411462 597134
rect 420226 597218 420462 597454
rect 420226 596898 420462 597134
rect 429226 597218 429462 597454
rect 429226 596898 429462 597134
rect 431788 597218 432024 597454
rect 431788 596898 432024 597134
rect 432440 597218 432676 597454
rect 432440 596898 432676 597134
rect 433246 597218 433482 597454
rect 433246 596898 433482 597134
rect 439792 597218 440028 597454
rect 439792 596898 440028 597134
rect 457010 597218 457246 597454
rect 457010 596898 457246 597134
rect 476652 597218 476888 597454
rect 476652 596898 476888 597134
rect 571716 597218 571952 597454
rect 571716 596898 571952 597134
rect 579470 597218 579706 597454
rect 579470 596898 579706 597134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect 5382 579218 5618 579454
rect 5382 578898 5618 579134
rect 13032 579218 13268 579454
rect 13032 578898 13268 579134
rect 106736 579218 106972 579454
rect 106736 578898 106972 579134
rect 127458 579218 127694 579454
rect 127458 578898 127694 579134
rect 140656 579218 140892 579454
rect 140656 578898 140892 579134
rect 141502 579218 141738 579454
rect 141502 578898 141738 579134
rect 147288 579218 147524 579454
rect 147288 578898 147524 579134
rect 149660 579218 149896 579454
rect 149660 578898 149896 579134
rect 150506 579218 150742 579454
rect 150506 578898 150742 579134
rect 159506 579218 159742 579454
rect 159506 578898 159742 579134
rect 168506 579218 168742 579454
rect 168506 578898 168742 579134
rect 177506 579218 177742 579454
rect 177506 578898 177742 579134
rect 186506 579218 186742 579454
rect 186506 578898 186742 579134
rect 188308 579218 188544 579454
rect 188308 578898 188544 579134
rect 190680 579218 190916 579454
rect 190680 578898 190916 579134
rect 191526 579218 191762 579454
rect 191526 578898 191762 579134
rect 200526 579218 200762 579454
rect 200526 578898 200762 579134
rect 209526 579218 209762 579454
rect 209526 578898 209762 579134
rect 218526 579218 218762 579454
rect 218526 578898 218762 579134
rect 227526 579218 227762 579454
rect 227526 578898 227762 579134
rect 229328 579218 229564 579454
rect 229328 578898 229564 579134
rect 230700 579218 230936 579454
rect 230700 578898 230936 579134
rect 231546 579218 231782 579454
rect 231546 578898 231782 579134
rect 240546 579218 240782 579454
rect 240546 578898 240782 579134
rect 249546 579218 249782 579454
rect 249546 578898 249782 579134
rect 258546 579218 258782 579454
rect 258546 578898 258782 579134
rect 267546 579218 267782 579454
rect 267546 578898 267782 579134
rect 269348 579218 269584 579454
rect 269348 578898 269584 579134
rect 270720 579218 270956 579454
rect 270720 578898 270956 579134
rect 271566 579218 271802 579454
rect 271566 578898 271802 579134
rect 280566 579218 280802 579454
rect 280566 578898 280802 579134
rect 289566 579218 289802 579454
rect 289566 578898 289802 579134
rect 298566 579218 298802 579454
rect 298566 578898 298802 579134
rect 307566 579218 307802 579454
rect 307566 578898 307802 579134
rect 309368 579218 309604 579454
rect 309368 578898 309604 579134
rect 311740 579218 311976 579454
rect 311740 578898 311976 579134
rect 312586 579218 312822 579454
rect 312586 578898 312822 579134
rect 321586 579218 321822 579454
rect 321586 578898 321822 579134
rect 330586 579218 330822 579454
rect 330586 578898 330822 579134
rect 339586 579218 339822 579454
rect 339586 578898 339822 579134
rect 348586 579218 348822 579454
rect 348586 578898 348822 579134
rect 350388 579218 350624 579454
rect 350388 578898 350624 579134
rect 352760 579218 352996 579454
rect 352760 578898 352996 579134
rect 353606 579218 353842 579454
rect 353606 578898 353842 579134
rect 362606 579218 362842 579454
rect 362606 578898 362842 579134
rect 371606 579218 371842 579454
rect 371606 578898 371842 579134
rect 380606 579218 380842 579454
rect 380606 578898 380842 579134
rect 389606 579218 389842 579454
rect 389606 578898 389842 579134
rect 391408 579218 391644 579454
rect 391408 578898 391644 579134
rect 392780 579218 393016 579454
rect 392780 578898 393016 579134
rect 393626 579218 393862 579454
rect 393626 578898 393862 579134
rect 402626 579218 402862 579454
rect 402626 578898 402862 579134
rect 411626 579218 411862 579454
rect 411626 578898 411862 579134
rect 420626 579218 420862 579454
rect 420626 578898 420862 579134
rect 429626 579218 429862 579454
rect 429626 578898 429862 579134
rect 431428 579218 431664 579454
rect 431428 578898 431664 579134
rect 432800 579218 433036 579454
rect 432800 578898 433036 579134
rect 433646 579218 433882 579454
rect 433646 578898 433882 579134
rect 439432 579218 439668 579454
rect 439432 578898 439668 579134
rect 456610 579218 456846 579454
rect 456610 578898 456846 579134
rect 477332 579218 477568 579454
rect 477332 578898 477568 579134
rect 571036 579218 571272 579454
rect 571036 578898 571272 579134
rect 578670 579218 578906 579454
rect 578670 578898 578906 579134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 4582 561218 4818 561454
rect 4582 560898 4818 561134
rect 12352 561218 12588 561454
rect 12352 560898 12588 561134
rect 107416 561218 107652 561454
rect 107416 560898 107652 561134
rect 127058 561218 127294 561454
rect 127058 560898 127294 561134
rect 140296 561218 140532 561454
rect 140296 560898 140532 561134
rect 141102 561218 141338 561454
rect 141102 560898 141338 561134
rect 147648 561218 147884 561454
rect 147648 560898 147884 561134
rect 149300 561218 149536 561454
rect 149300 560898 149536 561134
rect 150106 561218 150342 561454
rect 150106 560898 150342 561134
rect 159106 561218 159342 561454
rect 159106 560898 159342 561134
rect 168106 561218 168342 561454
rect 168106 560898 168342 561134
rect 177106 561218 177342 561454
rect 177106 560898 177342 561134
rect 186106 561218 186342 561454
rect 186106 560898 186342 561134
rect 188668 561218 188904 561454
rect 188668 560898 188904 561134
rect 190320 561218 190556 561454
rect 190320 560898 190556 561134
rect 191126 561218 191362 561454
rect 191126 560898 191362 561134
rect 200126 561218 200362 561454
rect 200126 560898 200362 561134
rect 209126 561218 209362 561454
rect 209126 560898 209362 561134
rect 218126 561218 218362 561454
rect 218126 560898 218362 561134
rect 227126 561218 227362 561454
rect 227126 560898 227362 561134
rect 229688 561218 229924 561454
rect 229688 560898 229924 561134
rect 230340 561218 230576 561454
rect 230340 560898 230576 561134
rect 231146 561218 231382 561454
rect 231146 560898 231382 561134
rect 240146 561218 240382 561454
rect 240146 560898 240382 561134
rect 249146 561218 249382 561454
rect 249146 560898 249382 561134
rect 258146 561218 258382 561454
rect 258146 560898 258382 561134
rect 267146 561218 267382 561454
rect 267146 560898 267382 561134
rect 269708 561218 269944 561454
rect 269708 560898 269944 561134
rect 270360 561218 270596 561454
rect 270360 560898 270596 561134
rect 271166 561218 271402 561454
rect 271166 560898 271402 561134
rect 280166 561218 280402 561454
rect 280166 560898 280402 561134
rect 289166 561218 289402 561454
rect 289166 560898 289402 561134
rect 298166 561218 298402 561454
rect 298166 560898 298402 561134
rect 307166 561218 307402 561454
rect 307166 560898 307402 561134
rect 309728 561218 309964 561454
rect 309728 560898 309964 561134
rect 311380 561218 311616 561454
rect 311380 560898 311616 561134
rect 312186 561218 312422 561454
rect 312186 560898 312422 561134
rect 321186 561218 321422 561454
rect 321186 560898 321422 561134
rect 330186 561218 330422 561454
rect 330186 560898 330422 561134
rect 339186 561218 339422 561454
rect 339186 560898 339422 561134
rect 348186 561218 348422 561454
rect 348186 560898 348422 561134
rect 350748 561218 350984 561454
rect 350748 560898 350984 561134
rect 352400 561218 352636 561454
rect 352400 560898 352636 561134
rect 353206 561218 353442 561454
rect 353206 560898 353442 561134
rect 362206 561218 362442 561454
rect 362206 560898 362442 561134
rect 371206 561218 371442 561454
rect 371206 560898 371442 561134
rect 380206 561218 380442 561454
rect 380206 560898 380442 561134
rect 389206 561218 389442 561454
rect 389206 560898 389442 561134
rect 391768 561218 392004 561454
rect 391768 560898 392004 561134
rect 392420 561218 392656 561454
rect 392420 560898 392656 561134
rect 393226 561218 393462 561454
rect 393226 560898 393462 561134
rect 402226 561218 402462 561454
rect 402226 560898 402462 561134
rect 411226 561218 411462 561454
rect 411226 560898 411462 561134
rect 420226 561218 420462 561454
rect 420226 560898 420462 561134
rect 429226 561218 429462 561454
rect 429226 560898 429462 561134
rect 431788 561218 432024 561454
rect 431788 560898 432024 561134
rect 432440 561218 432676 561454
rect 432440 560898 432676 561134
rect 433246 561218 433482 561454
rect 433246 560898 433482 561134
rect 439792 561218 440028 561454
rect 439792 560898 440028 561134
rect 457010 561218 457246 561454
rect 457010 560898 457246 561134
rect 476652 561218 476888 561454
rect 476652 560898 476888 561134
rect 571716 561218 571952 561454
rect 571716 560898 571952 561134
rect 579470 561218 579706 561454
rect 579470 560898 579706 561134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect 5382 543218 5618 543454
rect 5382 542898 5618 543134
rect 127458 543218 127694 543454
rect 127458 542898 127694 543134
rect 140656 543218 140892 543454
rect 140656 542898 140892 543134
rect 141502 543218 141738 543454
rect 141502 542898 141738 543134
rect 147288 543218 147524 543454
rect 147288 542898 147524 543134
rect 149660 543218 149896 543454
rect 149660 542898 149896 543134
rect 150506 543218 150742 543454
rect 150506 542898 150742 543134
rect 159506 543218 159742 543454
rect 159506 542898 159742 543134
rect 168506 543218 168742 543454
rect 168506 542898 168742 543134
rect 177506 543218 177742 543454
rect 177506 542898 177742 543134
rect 186506 543218 186742 543454
rect 186506 542898 186742 543134
rect 188308 543218 188544 543454
rect 188308 542898 188544 543134
rect 190680 543218 190916 543454
rect 190680 542898 190916 543134
rect 191526 543218 191762 543454
rect 191526 542898 191762 543134
rect 200526 543218 200762 543454
rect 200526 542898 200762 543134
rect 209526 543218 209762 543454
rect 209526 542898 209762 543134
rect 218526 543218 218762 543454
rect 218526 542898 218762 543134
rect 227526 543218 227762 543454
rect 227526 542898 227762 543134
rect 229328 543218 229564 543454
rect 229328 542898 229564 543134
rect 230700 543218 230936 543454
rect 230700 542898 230936 543134
rect 231546 543218 231782 543454
rect 231546 542898 231782 543134
rect 240546 543218 240782 543454
rect 240546 542898 240782 543134
rect 249546 543218 249782 543454
rect 249546 542898 249782 543134
rect 258546 543218 258782 543454
rect 258546 542898 258782 543134
rect 267546 543218 267782 543454
rect 267546 542898 267782 543134
rect 269348 543218 269584 543454
rect 269348 542898 269584 543134
rect 270720 543218 270956 543454
rect 270720 542898 270956 543134
rect 271566 543218 271802 543454
rect 271566 542898 271802 543134
rect 280566 543218 280802 543454
rect 280566 542898 280802 543134
rect 289566 543218 289802 543454
rect 289566 542898 289802 543134
rect 298566 543218 298802 543454
rect 298566 542898 298802 543134
rect 307566 543218 307802 543454
rect 307566 542898 307802 543134
rect 309368 543218 309604 543454
rect 309368 542898 309604 543134
rect 311740 543218 311976 543454
rect 311740 542898 311976 543134
rect 312586 543218 312822 543454
rect 312586 542898 312822 543134
rect 321586 543218 321822 543454
rect 321586 542898 321822 543134
rect 330586 543218 330822 543454
rect 330586 542898 330822 543134
rect 339586 543218 339822 543454
rect 339586 542898 339822 543134
rect 348586 543218 348822 543454
rect 348586 542898 348822 543134
rect 350388 543218 350624 543454
rect 350388 542898 350624 543134
rect 352760 543218 352996 543454
rect 352760 542898 352996 543134
rect 353606 543218 353842 543454
rect 353606 542898 353842 543134
rect 362606 543218 362842 543454
rect 362606 542898 362842 543134
rect 371606 543218 371842 543454
rect 371606 542898 371842 543134
rect 380606 543218 380842 543454
rect 380606 542898 380842 543134
rect 389606 543218 389842 543454
rect 389606 542898 389842 543134
rect 391408 543218 391644 543454
rect 391408 542898 391644 543134
rect 392780 543218 393016 543454
rect 392780 542898 393016 543134
rect 393626 543218 393862 543454
rect 393626 542898 393862 543134
rect 402626 543218 402862 543454
rect 402626 542898 402862 543134
rect 411626 543218 411862 543454
rect 411626 542898 411862 543134
rect 420626 543218 420862 543454
rect 420626 542898 420862 543134
rect 429626 543218 429862 543454
rect 429626 542898 429862 543134
rect 431428 543218 431664 543454
rect 431428 542898 431664 543134
rect 432800 543218 433036 543454
rect 432800 542898 433036 543134
rect 433646 543218 433882 543454
rect 433646 542898 433882 543134
rect 439432 543218 439668 543454
rect 439432 542898 439668 543134
rect 456610 543218 456846 543454
rect 456610 542898 456846 543134
rect 578670 543218 578906 543454
rect 578670 542898 578906 543134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 4582 525218 4818 525454
rect 4582 524898 4818 525134
rect 127058 525218 127294 525454
rect 127058 524898 127294 525134
rect 140296 525218 140532 525454
rect 140296 524898 140532 525134
rect 141102 525218 141338 525454
rect 141102 524898 141338 525134
rect 147648 525218 147884 525454
rect 147648 524898 147884 525134
rect 149300 525218 149536 525454
rect 149300 524898 149536 525134
rect 150106 525218 150342 525454
rect 150106 524898 150342 525134
rect 159106 525218 159342 525454
rect 159106 524898 159342 525134
rect 168106 525218 168342 525454
rect 168106 524898 168342 525134
rect 177106 525218 177342 525454
rect 177106 524898 177342 525134
rect 186106 525218 186342 525454
rect 186106 524898 186342 525134
rect 188668 525218 188904 525454
rect 188668 524898 188904 525134
rect 190320 525218 190556 525454
rect 190320 524898 190556 525134
rect 191126 525218 191362 525454
rect 191126 524898 191362 525134
rect 200126 525218 200362 525454
rect 200126 524898 200362 525134
rect 209126 525218 209362 525454
rect 209126 524898 209362 525134
rect 218126 525218 218362 525454
rect 218126 524898 218362 525134
rect 227126 525218 227362 525454
rect 227126 524898 227362 525134
rect 229688 525218 229924 525454
rect 229688 524898 229924 525134
rect 230340 525218 230576 525454
rect 230340 524898 230576 525134
rect 231146 525218 231382 525454
rect 231146 524898 231382 525134
rect 240146 525218 240382 525454
rect 240146 524898 240382 525134
rect 249146 525218 249382 525454
rect 249146 524898 249382 525134
rect 258146 525218 258382 525454
rect 258146 524898 258382 525134
rect 267146 525218 267382 525454
rect 267146 524898 267382 525134
rect 269708 525218 269944 525454
rect 269708 524898 269944 525134
rect 270360 525218 270596 525454
rect 270360 524898 270596 525134
rect 271166 525218 271402 525454
rect 271166 524898 271402 525134
rect 280166 525218 280402 525454
rect 280166 524898 280402 525134
rect 289166 525218 289402 525454
rect 289166 524898 289402 525134
rect 298166 525218 298402 525454
rect 298166 524898 298402 525134
rect 307166 525218 307402 525454
rect 307166 524898 307402 525134
rect 309728 525218 309964 525454
rect 309728 524898 309964 525134
rect 311380 525218 311616 525454
rect 311380 524898 311616 525134
rect 312186 525218 312422 525454
rect 312186 524898 312422 525134
rect 321186 525218 321422 525454
rect 321186 524898 321422 525134
rect 330186 525218 330422 525454
rect 330186 524898 330422 525134
rect 339186 525218 339422 525454
rect 339186 524898 339422 525134
rect 348186 525218 348422 525454
rect 348186 524898 348422 525134
rect 350748 525218 350984 525454
rect 350748 524898 350984 525134
rect 352400 525218 352636 525454
rect 352400 524898 352636 525134
rect 353206 525218 353442 525454
rect 353206 524898 353442 525134
rect 362206 525218 362442 525454
rect 362206 524898 362442 525134
rect 371206 525218 371442 525454
rect 371206 524898 371442 525134
rect 380206 525218 380442 525454
rect 380206 524898 380442 525134
rect 389206 525218 389442 525454
rect 389206 524898 389442 525134
rect 391768 525218 392004 525454
rect 391768 524898 392004 525134
rect 392420 525218 392656 525454
rect 392420 524898 392656 525134
rect 393226 525218 393462 525454
rect 393226 524898 393462 525134
rect 402226 525218 402462 525454
rect 402226 524898 402462 525134
rect 411226 525218 411462 525454
rect 411226 524898 411462 525134
rect 420226 525218 420462 525454
rect 420226 524898 420462 525134
rect 429226 525218 429462 525454
rect 429226 524898 429462 525134
rect 431788 525218 432024 525454
rect 431788 524898 432024 525134
rect 432440 525218 432676 525454
rect 432440 524898 432676 525134
rect 433246 525218 433482 525454
rect 433246 524898 433482 525134
rect 439792 525218 440028 525454
rect 439792 524898 440028 525134
rect 457010 525218 457246 525454
rect 457010 524898 457246 525134
rect 579470 525218 579706 525454
rect 579470 524898 579706 525134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect 5382 507218 5618 507454
rect 5382 506898 5618 507134
rect 127458 507218 127694 507454
rect 127458 506898 127694 507134
rect 140656 507218 140892 507454
rect 140656 506898 140892 507134
rect 141502 507218 141738 507454
rect 141502 506898 141738 507134
rect 147288 507218 147524 507454
rect 147288 506898 147524 507134
rect 149660 507218 149896 507454
rect 149660 506898 149896 507134
rect 150506 507218 150742 507454
rect 150506 506898 150742 507134
rect 159506 507218 159742 507454
rect 159506 506898 159742 507134
rect 168506 507218 168742 507454
rect 168506 506898 168742 507134
rect 177506 507218 177742 507454
rect 177506 506898 177742 507134
rect 186506 507218 186742 507454
rect 186506 506898 186742 507134
rect 188308 507218 188544 507454
rect 188308 506898 188544 507134
rect 190680 507218 190916 507454
rect 190680 506898 190916 507134
rect 191526 507218 191762 507454
rect 191526 506898 191762 507134
rect 200526 507218 200762 507454
rect 200526 506898 200762 507134
rect 209526 507218 209762 507454
rect 209526 506898 209762 507134
rect 218526 507218 218762 507454
rect 218526 506898 218762 507134
rect 227526 507218 227762 507454
rect 227526 506898 227762 507134
rect 229328 507218 229564 507454
rect 229328 506898 229564 507134
rect 230700 507218 230936 507454
rect 230700 506898 230936 507134
rect 231546 507218 231782 507454
rect 231546 506898 231782 507134
rect 240546 507218 240782 507454
rect 240546 506898 240782 507134
rect 249546 507218 249782 507454
rect 249546 506898 249782 507134
rect 258546 507218 258782 507454
rect 258546 506898 258782 507134
rect 267546 507218 267782 507454
rect 267546 506898 267782 507134
rect 269348 507218 269584 507454
rect 269348 506898 269584 507134
rect 270720 507218 270956 507454
rect 270720 506898 270956 507134
rect 271566 507218 271802 507454
rect 271566 506898 271802 507134
rect 280566 507218 280802 507454
rect 280566 506898 280802 507134
rect 289566 507218 289802 507454
rect 289566 506898 289802 507134
rect 298566 507218 298802 507454
rect 298566 506898 298802 507134
rect 307566 507218 307802 507454
rect 307566 506898 307802 507134
rect 309368 507218 309604 507454
rect 309368 506898 309604 507134
rect 311740 507218 311976 507454
rect 311740 506898 311976 507134
rect 312586 507218 312822 507454
rect 312586 506898 312822 507134
rect 321586 507218 321822 507454
rect 321586 506898 321822 507134
rect 330586 507218 330822 507454
rect 330586 506898 330822 507134
rect 339586 507218 339822 507454
rect 339586 506898 339822 507134
rect 348586 507218 348822 507454
rect 348586 506898 348822 507134
rect 350388 507218 350624 507454
rect 350388 506898 350624 507134
rect 352760 507218 352996 507454
rect 352760 506898 352996 507134
rect 353606 507218 353842 507454
rect 353606 506898 353842 507134
rect 362606 507218 362842 507454
rect 362606 506898 362842 507134
rect 371606 507218 371842 507454
rect 371606 506898 371842 507134
rect 380606 507218 380842 507454
rect 380606 506898 380842 507134
rect 389606 507218 389842 507454
rect 389606 506898 389842 507134
rect 391408 507218 391644 507454
rect 391408 506898 391644 507134
rect 392780 507218 393016 507454
rect 392780 506898 393016 507134
rect 393626 507218 393862 507454
rect 393626 506898 393862 507134
rect 402626 507218 402862 507454
rect 402626 506898 402862 507134
rect 411626 507218 411862 507454
rect 411626 506898 411862 507134
rect 420626 507218 420862 507454
rect 420626 506898 420862 507134
rect 429626 507218 429862 507454
rect 429626 506898 429862 507134
rect 431428 507218 431664 507454
rect 431428 506898 431664 507134
rect 432800 507218 433036 507454
rect 432800 506898 433036 507134
rect 433646 507218 433882 507454
rect 433646 506898 433882 507134
rect 439432 507218 439668 507454
rect 439432 506898 439668 507134
rect 456610 507218 456846 507454
rect 456610 506898 456846 507134
rect 578670 507218 578906 507454
rect 578670 506898 578906 507134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 4582 489218 4818 489454
rect 4582 488898 4818 489134
rect 12618 489218 12854 489454
rect 12618 488898 12854 489134
rect 14040 489218 14276 489454
rect 14040 488898 14276 489134
rect 23040 489218 23276 489454
rect 23040 488898 23276 489134
rect 32040 489218 32276 489454
rect 32040 488898 32276 489134
rect 41040 489218 41276 489454
rect 41040 488898 41276 489134
rect 50040 489218 50276 489454
rect 50040 488898 50276 489134
rect 59040 489218 59276 489454
rect 59040 488898 59276 489134
rect 68040 489218 68276 489454
rect 68040 488898 68276 489134
rect 77040 489218 77276 489454
rect 77040 488898 77276 489134
rect 86040 489218 86276 489454
rect 86040 488898 86276 489134
rect 95040 489218 95276 489454
rect 95040 488898 95276 489134
rect 104040 489218 104276 489454
rect 104040 488898 104276 489134
rect 113040 489218 113276 489454
rect 113040 488898 113276 489134
rect 121226 489218 121462 489454
rect 121226 488898 121462 489134
rect 127058 489218 127294 489454
rect 127058 488898 127294 489134
rect 140296 489218 140532 489454
rect 140296 488898 140532 489134
rect 141102 489218 141338 489454
rect 141102 488898 141338 489134
rect 147648 489218 147884 489454
rect 147648 488898 147884 489134
rect 149300 489218 149536 489454
rect 149300 488898 149536 489134
rect 150106 489218 150342 489454
rect 150106 488898 150342 489134
rect 159106 489218 159342 489454
rect 159106 488898 159342 489134
rect 168106 489218 168342 489454
rect 168106 488898 168342 489134
rect 177106 489218 177342 489454
rect 177106 488898 177342 489134
rect 186106 489218 186342 489454
rect 186106 488898 186342 489134
rect 188668 489218 188904 489454
rect 188668 488898 188904 489134
rect 189768 489218 190004 489454
rect 189768 488898 190004 489134
rect 190320 489218 190556 489454
rect 190320 488898 190556 489134
rect 191126 489218 191362 489454
rect 191126 488898 191362 489134
rect 200126 489218 200362 489454
rect 200126 488898 200362 489134
rect 209126 489218 209362 489454
rect 209126 488898 209362 489134
rect 218126 489218 218362 489454
rect 218126 488898 218362 489134
rect 227126 489218 227362 489454
rect 227126 488898 227362 489134
rect 229688 489218 229924 489454
rect 229688 488898 229924 489134
rect 230340 489218 230576 489454
rect 230340 488898 230576 489134
rect 231146 489218 231382 489454
rect 231146 488898 231382 489134
rect 240146 489218 240382 489454
rect 240146 488898 240382 489134
rect 249146 489218 249382 489454
rect 249146 488898 249382 489134
rect 258146 489218 258382 489454
rect 258146 488898 258382 489134
rect 267146 489218 267382 489454
rect 267146 488898 267382 489134
rect 269708 489218 269944 489454
rect 269708 488898 269944 489134
rect 270360 489218 270596 489454
rect 270360 488898 270596 489134
rect 271166 489218 271402 489454
rect 271166 488898 271402 489134
rect 280166 489218 280402 489454
rect 280166 488898 280402 489134
rect 289166 489218 289402 489454
rect 289166 488898 289402 489134
rect 298166 489218 298402 489454
rect 298166 488898 298402 489134
rect 307166 489218 307402 489454
rect 307166 488898 307402 489134
rect 309728 489218 309964 489454
rect 309728 488898 309964 489134
rect 311380 489218 311616 489454
rect 311380 488898 311616 489134
rect 312186 489218 312422 489454
rect 312186 488898 312422 489134
rect 321186 489218 321422 489454
rect 321186 488898 321422 489134
rect 330186 489218 330422 489454
rect 330186 488898 330422 489134
rect 339186 489218 339422 489454
rect 339186 488898 339422 489134
rect 348186 489218 348422 489454
rect 348186 488898 348422 489134
rect 350748 489218 350984 489454
rect 350748 488898 350984 489134
rect 352400 489218 352636 489454
rect 352400 488898 352636 489134
rect 353206 489218 353442 489454
rect 353206 488898 353442 489134
rect 362206 489218 362442 489454
rect 362206 488898 362442 489134
rect 371206 489218 371442 489454
rect 371206 488898 371442 489134
rect 380206 489218 380442 489454
rect 380206 488898 380442 489134
rect 389206 489218 389442 489454
rect 389206 488898 389442 489134
rect 391768 489218 392004 489454
rect 391768 488898 392004 489134
rect 392420 489218 392656 489454
rect 392420 488898 392656 489134
rect 393226 489218 393462 489454
rect 393226 488898 393462 489134
rect 402226 489218 402462 489454
rect 402226 488898 402462 489134
rect 411226 489218 411462 489454
rect 411226 488898 411462 489134
rect 420226 489218 420462 489454
rect 420226 488898 420462 489134
rect 429226 489218 429462 489454
rect 429226 488898 429462 489134
rect 431788 489218 432024 489454
rect 431788 488898 432024 489134
rect 432440 489218 432676 489454
rect 432440 488898 432676 489134
rect 433246 489218 433482 489454
rect 433246 488898 433482 489134
rect 439792 489218 440028 489454
rect 439792 488898 440028 489134
rect 457010 489218 457246 489454
rect 457010 488898 457246 489134
rect 462842 489218 463078 489454
rect 462842 488898 463078 489134
rect 471028 489218 471264 489454
rect 471028 488898 471264 489134
rect 480028 489218 480264 489454
rect 480028 488898 480264 489134
rect 489028 489218 489264 489454
rect 489028 488898 489264 489134
rect 498028 489218 498264 489454
rect 498028 488898 498264 489134
rect 507028 489218 507264 489454
rect 507028 488898 507264 489134
rect 516028 489218 516264 489454
rect 516028 488898 516264 489134
rect 525028 489218 525264 489454
rect 525028 488898 525264 489134
rect 534028 489218 534264 489454
rect 534028 488898 534264 489134
rect 543028 489218 543264 489454
rect 543028 488898 543264 489134
rect 552028 489218 552264 489454
rect 552028 488898 552264 489134
rect 561028 489218 561264 489454
rect 561028 488898 561264 489134
rect 570028 489218 570264 489454
rect 570028 488898 570264 489134
rect 571450 489218 571686 489454
rect 571450 488898 571686 489134
rect 579470 489218 579706 489454
rect 579470 488898 579706 489134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect 5382 471218 5618 471454
rect 5382 470898 5618 471134
rect 13218 471218 13454 471454
rect 13218 470898 13454 471134
rect 14420 471218 14656 471454
rect 14420 470898 14656 471134
rect 23420 471218 23656 471454
rect 23420 470898 23656 471134
rect 32420 471218 32656 471454
rect 32420 470898 32656 471134
rect 41420 471218 41656 471454
rect 41420 470898 41656 471134
rect 50420 471218 50656 471454
rect 50420 470898 50656 471134
rect 59420 471218 59656 471454
rect 59420 470898 59656 471134
rect 68420 471218 68656 471454
rect 68420 470898 68656 471134
rect 77420 471218 77656 471454
rect 77420 470898 77656 471134
rect 86420 471218 86656 471454
rect 86420 470898 86656 471134
rect 95420 471218 95656 471454
rect 95420 470898 95656 471134
rect 104420 471218 104656 471454
rect 104420 470898 104656 471134
rect 113420 471218 113656 471454
rect 113420 470898 113656 471134
rect 120626 471218 120862 471454
rect 120626 470898 120862 471134
rect 127458 471218 127694 471454
rect 127458 470898 127694 471134
rect 140656 471218 140892 471454
rect 140656 470898 140892 471134
rect 141502 471218 141738 471454
rect 141502 470898 141738 471134
rect 147288 471218 147524 471454
rect 147288 470898 147524 471134
rect 149660 471218 149896 471454
rect 149660 470898 149896 471134
rect 150506 471218 150742 471454
rect 150506 470898 150742 471134
rect 159506 471218 159742 471454
rect 159506 470898 159742 471134
rect 168506 471218 168742 471454
rect 168506 470898 168742 471134
rect 177506 471218 177742 471454
rect 177506 470898 177742 471134
rect 186506 471218 186742 471454
rect 186506 470898 186742 471134
rect 188308 471218 188544 471454
rect 188308 470898 188544 471134
rect 190680 471218 190916 471454
rect 190680 470898 190916 471134
rect 191526 471218 191762 471454
rect 191526 470898 191762 471134
rect 200526 471218 200762 471454
rect 200526 470898 200762 471134
rect 209526 471218 209762 471454
rect 209526 470898 209762 471134
rect 218526 471218 218762 471454
rect 218526 470898 218762 471134
rect 227526 471218 227762 471454
rect 227526 470898 227762 471134
rect 229328 471218 229564 471454
rect 229328 470898 229564 471134
rect 230700 471218 230936 471454
rect 230700 470898 230936 471134
rect 231546 471218 231782 471454
rect 231546 470898 231782 471134
rect 240546 471218 240782 471454
rect 240546 470898 240782 471134
rect 249546 471218 249782 471454
rect 249546 470898 249782 471134
rect 258546 471218 258782 471454
rect 258546 470898 258782 471134
rect 267546 471218 267782 471454
rect 267546 470898 267782 471134
rect 269348 471218 269584 471454
rect 269348 470898 269584 471134
rect 270720 471218 270956 471454
rect 270720 470898 270956 471134
rect 271566 471218 271802 471454
rect 271566 470898 271802 471134
rect 280566 471218 280802 471454
rect 280566 470898 280802 471134
rect 289566 471218 289802 471454
rect 289566 470898 289802 471134
rect 298566 471218 298802 471454
rect 298566 470898 298802 471134
rect 307566 471218 307802 471454
rect 307566 470898 307802 471134
rect 309368 471218 309604 471454
rect 309368 470898 309604 471134
rect 311740 471218 311976 471454
rect 311740 470898 311976 471134
rect 312586 471218 312822 471454
rect 312586 470898 312822 471134
rect 321586 471218 321822 471454
rect 321586 470898 321822 471134
rect 330586 471218 330822 471454
rect 330586 470898 330822 471134
rect 339586 471218 339822 471454
rect 339586 470898 339822 471134
rect 348586 471218 348822 471454
rect 348586 470898 348822 471134
rect 350388 471218 350624 471454
rect 350388 470898 350624 471134
rect 352760 471218 352996 471454
rect 352760 470898 352996 471134
rect 353606 471218 353842 471454
rect 353606 470898 353842 471134
rect 362606 471218 362842 471454
rect 362606 470898 362842 471134
rect 371606 471218 371842 471454
rect 371606 470898 371842 471134
rect 380606 471218 380842 471454
rect 380606 470898 380842 471134
rect 389606 471218 389842 471454
rect 389606 470898 389842 471134
rect 391408 471218 391644 471454
rect 391408 470898 391644 471134
rect 392780 471218 393016 471454
rect 392780 470898 393016 471134
rect 393626 471218 393862 471454
rect 393626 470898 393862 471134
rect 402626 471218 402862 471454
rect 402626 470898 402862 471134
rect 411626 471218 411862 471454
rect 411626 470898 411862 471134
rect 420626 471218 420862 471454
rect 420626 470898 420862 471134
rect 429626 471218 429862 471454
rect 429626 470898 429862 471134
rect 431428 471218 431664 471454
rect 431428 470898 431664 471134
rect 432800 471218 433036 471454
rect 432800 470898 433036 471134
rect 433646 471218 433882 471454
rect 433646 470898 433882 471134
rect 439432 471218 439668 471454
rect 439432 470898 439668 471134
rect 456610 471218 456846 471454
rect 456610 470898 456846 471134
rect 463442 471218 463678 471454
rect 463442 470898 463678 471134
rect 470648 471218 470884 471454
rect 470648 470898 470884 471134
rect 479648 471218 479884 471454
rect 479648 470898 479884 471134
rect 488648 471218 488884 471454
rect 488648 470898 488884 471134
rect 497648 471218 497884 471454
rect 497648 470898 497884 471134
rect 506648 471218 506884 471454
rect 506648 470898 506884 471134
rect 515648 471218 515884 471454
rect 515648 470898 515884 471134
rect 524648 471218 524884 471454
rect 524648 470898 524884 471134
rect 533648 471218 533884 471454
rect 533648 470898 533884 471134
rect 542648 471218 542884 471454
rect 542648 470898 542884 471134
rect 551648 471218 551884 471454
rect 551648 470898 551884 471134
rect 560648 471218 560884 471454
rect 560648 470898 560884 471134
rect 569648 471218 569884 471454
rect 569648 470898 569884 471134
rect 570850 471218 571086 471454
rect 570850 470898 571086 471134
rect 578670 471218 578906 471454
rect 578670 470898 578906 471134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 4582 453218 4818 453454
rect 4582 452898 4818 453134
rect 12618 453218 12854 453454
rect 12618 452898 12854 453134
rect 14040 453218 14276 453454
rect 14040 452898 14276 453134
rect 23040 453218 23276 453454
rect 23040 452898 23276 453134
rect 32040 453218 32276 453454
rect 32040 452898 32276 453134
rect 41040 453218 41276 453454
rect 41040 452898 41276 453134
rect 50040 453218 50276 453454
rect 50040 452898 50276 453134
rect 59040 453218 59276 453454
rect 59040 452898 59276 453134
rect 68040 453218 68276 453454
rect 68040 452898 68276 453134
rect 77040 453218 77276 453454
rect 77040 452898 77276 453134
rect 86040 453218 86276 453454
rect 86040 452898 86276 453134
rect 95040 453218 95276 453454
rect 95040 452898 95276 453134
rect 104040 453218 104276 453454
rect 104040 452898 104276 453134
rect 113040 453218 113276 453454
rect 113040 452898 113276 453134
rect 121226 453218 121462 453454
rect 121226 452898 121462 453134
rect 127058 453218 127294 453454
rect 127058 452898 127294 453134
rect 140296 453218 140532 453454
rect 140296 452898 140532 453134
rect 141102 453218 141338 453454
rect 141102 452898 141338 453134
rect 147648 453218 147884 453454
rect 147648 452898 147884 453134
rect 149300 453218 149536 453454
rect 149300 452898 149536 453134
rect 150106 453218 150342 453454
rect 150106 452898 150342 453134
rect 159106 453218 159342 453454
rect 159106 452898 159342 453134
rect 168106 453218 168342 453454
rect 168106 452898 168342 453134
rect 177106 453218 177342 453454
rect 177106 452898 177342 453134
rect 186106 453218 186342 453454
rect 186106 452898 186342 453134
rect 188668 453218 188904 453454
rect 188668 452898 188904 453134
rect 190320 453218 190556 453454
rect 190320 452898 190556 453134
rect 191126 453218 191362 453454
rect 191126 452898 191362 453134
rect 200126 453218 200362 453454
rect 200126 452898 200362 453134
rect 209126 453218 209362 453454
rect 209126 452898 209362 453134
rect 218126 453218 218362 453454
rect 218126 452898 218362 453134
rect 227126 453218 227362 453454
rect 227126 452898 227362 453134
rect 229688 453218 229924 453454
rect 229688 452898 229924 453134
rect 230340 453218 230576 453454
rect 230340 452898 230576 453134
rect 231146 453218 231382 453454
rect 231146 452898 231382 453134
rect 240146 453218 240382 453454
rect 240146 452898 240382 453134
rect 249146 453218 249382 453454
rect 249146 452898 249382 453134
rect 258146 453218 258382 453454
rect 258146 452898 258382 453134
rect 267146 453218 267382 453454
rect 267146 452898 267382 453134
rect 269708 453218 269944 453454
rect 269708 452898 269944 453134
rect 270360 453218 270596 453454
rect 270360 452898 270596 453134
rect 271166 453218 271402 453454
rect 271166 452898 271402 453134
rect 280166 453218 280402 453454
rect 280166 452898 280402 453134
rect 289166 453218 289402 453454
rect 289166 452898 289402 453134
rect 298166 453218 298402 453454
rect 298166 452898 298402 453134
rect 307166 453218 307402 453454
rect 307166 452898 307402 453134
rect 309728 453218 309964 453454
rect 309728 452898 309964 453134
rect 311380 453218 311616 453454
rect 311380 452898 311616 453134
rect 312186 453218 312422 453454
rect 312186 452898 312422 453134
rect 321186 453218 321422 453454
rect 321186 452898 321422 453134
rect 330186 453218 330422 453454
rect 330186 452898 330422 453134
rect 339186 453218 339422 453454
rect 339186 452898 339422 453134
rect 348186 453218 348422 453454
rect 348186 452898 348422 453134
rect 350748 453218 350984 453454
rect 350748 452898 350984 453134
rect 352400 453218 352636 453454
rect 352400 452898 352636 453134
rect 353206 453218 353442 453454
rect 353206 452898 353442 453134
rect 362206 453218 362442 453454
rect 362206 452898 362442 453134
rect 371206 453218 371442 453454
rect 371206 452898 371442 453134
rect 380206 453218 380442 453454
rect 380206 452898 380442 453134
rect 389206 453218 389442 453454
rect 389206 452898 389442 453134
rect 391768 453218 392004 453454
rect 391768 452898 392004 453134
rect 392420 453218 392656 453454
rect 392420 452898 392656 453134
rect 393226 453218 393462 453454
rect 393226 452898 393462 453134
rect 402226 453218 402462 453454
rect 402226 452898 402462 453134
rect 411226 453218 411462 453454
rect 411226 452898 411462 453134
rect 420226 453218 420462 453454
rect 420226 452898 420462 453134
rect 429226 453218 429462 453454
rect 429226 452898 429462 453134
rect 431788 453218 432024 453454
rect 431788 452898 432024 453134
rect 432440 453218 432676 453454
rect 432440 452898 432676 453134
rect 433246 453218 433482 453454
rect 433246 452898 433482 453134
rect 439792 453218 440028 453454
rect 439792 452898 440028 453134
rect 457010 453218 457246 453454
rect 457010 452898 457246 453134
rect 462842 453218 463078 453454
rect 462842 452898 463078 453134
rect 471028 453218 471264 453454
rect 471028 452898 471264 453134
rect 480028 453218 480264 453454
rect 480028 452898 480264 453134
rect 489028 453218 489264 453454
rect 489028 452898 489264 453134
rect 498028 453218 498264 453454
rect 498028 452898 498264 453134
rect 507028 453218 507264 453454
rect 507028 452898 507264 453134
rect 516028 453218 516264 453454
rect 516028 452898 516264 453134
rect 525028 453218 525264 453454
rect 525028 452898 525264 453134
rect 534028 453218 534264 453454
rect 534028 452898 534264 453134
rect 543028 453218 543264 453454
rect 543028 452898 543264 453134
rect 552028 453218 552264 453454
rect 552028 452898 552264 453134
rect 561028 453218 561264 453454
rect 561028 452898 561264 453134
rect 570028 453218 570264 453454
rect 570028 452898 570264 453134
rect 571450 453218 571686 453454
rect 571450 452898 571686 453134
rect 579470 453218 579706 453454
rect 579470 452898 579706 453134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect 5382 435218 5618 435454
rect 5382 434898 5618 435134
rect 13218 435218 13454 435454
rect 13218 434898 13454 435134
rect 14420 435218 14656 435454
rect 14420 434898 14656 435134
rect 23420 435218 23656 435454
rect 23420 434898 23656 435134
rect 32420 435218 32656 435454
rect 32420 434898 32656 435134
rect 41420 435218 41656 435454
rect 41420 434898 41656 435134
rect 50420 435218 50656 435454
rect 50420 434898 50656 435134
rect 59420 435218 59656 435454
rect 59420 434898 59656 435134
rect 68420 435218 68656 435454
rect 68420 434898 68656 435134
rect 77420 435218 77656 435454
rect 77420 434898 77656 435134
rect 86420 435218 86656 435454
rect 86420 434898 86656 435134
rect 95420 435218 95656 435454
rect 95420 434898 95656 435134
rect 104420 435218 104656 435454
rect 104420 434898 104656 435134
rect 113420 435218 113656 435454
rect 113420 434898 113656 435134
rect 120626 435218 120862 435454
rect 120626 434898 120862 435134
rect 127458 435218 127694 435454
rect 127458 434898 127694 435134
rect 140656 435218 140892 435454
rect 140656 434898 140892 435134
rect 147288 435218 147524 435454
rect 147288 434898 147524 435134
rect 149660 435218 149896 435454
rect 149660 434898 149896 435134
rect 150506 435218 150742 435454
rect 150506 434898 150742 435134
rect 159506 435218 159742 435454
rect 159506 434898 159742 435134
rect 168506 435218 168742 435454
rect 168506 434898 168742 435134
rect 177506 435218 177742 435454
rect 177506 434898 177742 435134
rect 186506 435218 186742 435454
rect 186506 434898 186742 435134
rect 188308 435218 188544 435454
rect 188308 434898 188544 435134
rect 190680 435218 190916 435454
rect 190680 434898 190916 435134
rect 229328 435218 229564 435454
rect 229328 434898 229564 435134
rect 230700 435218 230936 435454
rect 230700 434898 230936 435134
rect 269348 435218 269584 435454
rect 269348 434898 269584 435134
rect 270720 435218 270956 435454
rect 270720 434898 270956 435134
rect 309368 435218 309604 435454
rect 309368 434898 309604 435134
rect 311740 435218 311976 435454
rect 311740 434898 311976 435134
rect 312586 435218 312822 435454
rect 312586 434898 312822 435134
rect 321586 435218 321822 435454
rect 321586 434898 321822 435134
rect 330586 435218 330822 435454
rect 330586 434898 330822 435134
rect 339586 435218 339822 435454
rect 339586 434898 339822 435134
rect 348586 435218 348822 435454
rect 348586 434898 348822 435134
rect 350388 435218 350624 435454
rect 350388 434898 350624 435134
rect 352760 435218 352996 435454
rect 352760 434898 352996 435134
rect 391408 435218 391644 435454
rect 391408 434898 391644 435134
rect 392780 435218 393016 435454
rect 392780 434898 393016 435134
rect 431428 435218 431664 435454
rect 431428 434898 431664 435134
rect 432800 435218 433036 435454
rect 432800 434898 433036 435134
rect 439432 435218 439668 435454
rect 439432 434898 439668 435134
rect 456610 435218 456846 435454
rect 456610 434898 456846 435134
rect 463442 435218 463678 435454
rect 463442 434898 463678 435134
rect 470648 435218 470884 435454
rect 470648 434898 470884 435134
rect 479648 435218 479884 435454
rect 479648 434898 479884 435134
rect 488648 435218 488884 435454
rect 488648 434898 488884 435134
rect 497648 435218 497884 435454
rect 497648 434898 497884 435134
rect 506648 435218 506884 435454
rect 506648 434898 506884 435134
rect 515648 435218 515884 435454
rect 515648 434898 515884 435134
rect 524648 435218 524884 435454
rect 524648 434898 524884 435134
rect 533648 435218 533884 435454
rect 533648 434898 533884 435134
rect 542648 435218 542884 435454
rect 542648 434898 542884 435134
rect 551648 435218 551884 435454
rect 551648 434898 551884 435134
rect 560648 435218 560884 435454
rect 560648 434898 560884 435134
rect 569648 435218 569884 435454
rect 569648 434898 569884 435134
rect 570850 435218 571086 435454
rect 570850 434898 571086 435134
rect 578670 435218 578906 435454
rect 578670 434898 578906 435134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 4582 417218 4818 417454
rect 4582 416898 4818 417134
rect 12618 417218 12854 417454
rect 12618 416898 12854 417134
rect 14040 417218 14276 417454
rect 14040 416898 14276 417134
rect 23040 417218 23276 417454
rect 23040 416898 23276 417134
rect 32040 417218 32276 417454
rect 32040 416898 32276 417134
rect 41040 417218 41276 417454
rect 41040 416898 41276 417134
rect 50040 417218 50276 417454
rect 50040 416898 50276 417134
rect 59040 417218 59276 417454
rect 59040 416898 59276 417134
rect 68040 417218 68276 417454
rect 68040 416898 68276 417134
rect 77040 417218 77276 417454
rect 77040 416898 77276 417134
rect 86040 417218 86276 417454
rect 86040 416898 86276 417134
rect 95040 417218 95276 417454
rect 95040 416898 95276 417134
rect 104040 417218 104276 417454
rect 104040 416898 104276 417134
rect 113040 417218 113276 417454
rect 113040 416898 113276 417134
rect 121226 417218 121462 417454
rect 121226 416898 121462 417134
rect 127058 417218 127294 417454
rect 127058 416898 127294 417134
rect 140296 417218 140532 417454
rect 140296 416898 140532 417134
rect 141102 417218 141338 417454
rect 141102 416898 141338 417134
rect 147648 417218 147884 417454
rect 147648 416898 147884 417134
rect 149300 417218 149536 417454
rect 149300 416898 149536 417134
rect 150106 417218 150342 417454
rect 150106 416898 150342 417134
rect 159106 417218 159342 417454
rect 159106 416898 159342 417134
rect 168106 417218 168342 417454
rect 168106 416898 168342 417134
rect 177106 417218 177342 417454
rect 177106 416898 177342 417134
rect 186106 417218 186342 417454
rect 186106 416898 186342 417134
rect 188668 417218 188904 417454
rect 188668 416898 188904 417134
rect 189768 417218 190004 417454
rect 189768 416898 190004 417134
rect 190320 417218 190556 417454
rect 190320 416898 190556 417134
rect 191126 417218 191362 417454
rect 191126 416898 191362 417134
rect 200126 417218 200362 417454
rect 200126 416898 200362 417134
rect 209126 417218 209362 417454
rect 209126 416898 209362 417134
rect 218126 417218 218362 417454
rect 218126 416898 218362 417134
rect 227126 417218 227362 417454
rect 227126 416898 227362 417134
rect 229688 417218 229924 417454
rect 229688 416898 229924 417134
rect 230340 417218 230576 417454
rect 230340 416898 230576 417134
rect 231146 417218 231382 417454
rect 231146 416898 231382 417134
rect 240146 417218 240382 417454
rect 240146 416898 240382 417134
rect 249146 417218 249382 417454
rect 249146 416898 249382 417134
rect 258146 417218 258382 417454
rect 258146 416898 258382 417134
rect 267146 417218 267382 417454
rect 267146 416898 267382 417134
rect 269708 417218 269944 417454
rect 269708 416898 269944 417134
rect 270360 417218 270596 417454
rect 270360 416898 270596 417134
rect 271166 417218 271402 417454
rect 271166 416898 271402 417134
rect 280166 417218 280402 417454
rect 280166 416898 280402 417134
rect 289166 417218 289402 417454
rect 289166 416898 289402 417134
rect 298166 417218 298402 417454
rect 298166 416898 298402 417134
rect 307166 417218 307402 417454
rect 307166 416898 307402 417134
rect 309728 417218 309964 417454
rect 309728 416898 309964 417134
rect 311380 417218 311616 417454
rect 311380 416898 311616 417134
rect 312186 417218 312422 417454
rect 312186 416898 312422 417134
rect 321186 417218 321422 417454
rect 321186 416898 321422 417134
rect 330186 417218 330422 417454
rect 330186 416898 330422 417134
rect 339186 417218 339422 417454
rect 339186 416898 339422 417134
rect 348186 417218 348422 417454
rect 348186 416898 348422 417134
rect 350748 417218 350984 417454
rect 350748 416898 350984 417134
rect 352400 417218 352636 417454
rect 352400 416898 352636 417134
rect 353206 417218 353442 417454
rect 353206 416898 353442 417134
rect 362206 417218 362442 417454
rect 362206 416898 362442 417134
rect 371206 417218 371442 417454
rect 371206 416898 371442 417134
rect 380206 417218 380442 417454
rect 380206 416898 380442 417134
rect 389206 417218 389442 417454
rect 389206 416898 389442 417134
rect 391768 417218 392004 417454
rect 391768 416898 392004 417134
rect 392420 417218 392656 417454
rect 392420 416898 392656 417134
rect 393226 417218 393462 417454
rect 393226 416898 393462 417134
rect 402226 417218 402462 417454
rect 402226 416898 402462 417134
rect 411226 417218 411462 417454
rect 411226 416898 411462 417134
rect 420226 417218 420462 417454
rect 420226 416898 420462 417134
rect 429226 417218 429462 417454
rect 429226 416898 429462 417134
rect 431788 417218 432024 417454
rect 431788 416898 432024 417134
rect 432440 417218 432676 417454
rect 432440 416898 432676 417134
rect 433246 417218 433482 417454
rect 433246 416898 433482 417134
rect 439792 417218 440028 417454
rect 439792 416898 440028 417134
rect 457010 417218 457246 417454
rect 457010 416898 457246 417134
rect 462842 417218 463078 417454
rect 462842 416898 463078 417134
rect 471028 417218 471264 417454
rect 471028 416898 471264 417134
rect 480028 417218 480264 417454
rect 480028 416898 480264 417134
rect 489028 417218 489264 417454
rect 489028 416898 489264 417134
rect 498028 417218 498264 417454
rect 498028 416898 498264 417134
rect 507028 417218 507264 417454
rect 507028 416898 507264 417134
rect 516028 417218 516264 417454
rect 516028 416898 516264 417134
rect 525028 417218 525264 417454
rect 525028 416898 525264 417134
rect 534028 417218 534264 417454
rect 534028 416898 534264 417134
rect 543028 417218 543264 417454
rect 543028 416898 543264 417134
rect 552028 417218 552264 417454
rect 552028 416898 552264 417134
rect 561028 417218 561264 417454
rect 561028 416898 561264 417134
rect 570028 417218 570264 417454
rect 570028 416898 570264 417134
rect 571450 417218 571686 417454
rect 571450 416898 571686 417134
rect 579470 417218 579706 417454
rect 579470 416898 579706 417134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect 5382 399218 5618 399454
rect 5382 398898 5618 399134
rect 13218 399218 13454 399454
rect 13218 398898 13454 399134
rect 14420 399218 14656 399454
rect 14420 398898 14656 399134
rect 23420 399218 23656 399454
rect 23420 398898 23656 399134
rect 32420 399218 32656 399454
rect 32420 398898 32656 399134
rect 41420 399218 41656 399454
rect 41420 398898 41656 399134
rect 50420 399218 50656 399454
rect 50420 398898 50656 399134
rect 59420 399218 59656 399454
rect 59420 398898 59656 399134
rect 68420 399218 68656 399454
rect 68420 398898 68656 399134
rect 77420 399218 77656 399454
rect 77420 398898 77656 399134
rect 86420 399218 86656 399454
rect 86420 398898 86656 399134
rect 95420 399218 95656 399454
rect 95420 398898 95656 399134
rect 104420 399218 104656 399454
rect 104420 398898 104656 399134
rect 113420 399218 113656 399454
rect 113420 398898 113656 399134
rect 120626 399218 120862 399454
rect 120626 398898 120862 399134
rect 127458 399218 127694 399454
rect 127458 398898 127694 399134
rect 140656 399218 140892 399454
rect 140656 398898 140892 399134
rect 141502 399218 141738 399454
rect 141502 398898 141738 399134
rect 147288 399218 147524 399454
rect 147288 398898 147524 399134
rect 149660 399218 149896 399454
rect 149660 398898 149896 399134
rect 150506 399218 150742 399454
rect 150506 398898 150742 399134
rect 159506 399218 159742 399454
rect 159506 398898 159742 399134
rect 168506 399218 168742 399454
rect 168506 398898 168742 399134
rect 177506 399218 177742 399454
rect 177506 398898 177742 399134
rect 186506 399218 186742 399454
rect 186506 398898 186742 399134
rect 188308 399218 188544 399454
rect 188308 398898 188544 399134
rect 190680 399218 190916 399454
rect 190680 398898 190916 399134
rect 191526 399218 191762 399454
rect 191526 398898 191762 399134
rect 200526 399218 200762 399454
rect 200526 398898 200762 399134
rect 209526 399218 209762 399454
rect 209526 398898 209762 399134
rect 218526 399218 218762 399454
rect 218526 398898 218762 399134
rect 227526 399218 227762 399454
rect 227526 398898 227762 399134
rect 229328 399218 229564 399454
rect 229328 398898 229564 399134
rect 230700 399218 230936 399454
rect 230700 398898 230936 399134
rect 231546 399218 231782 399454
rect 231546 398898 231782 399134
rect 240546 399218 240782 399454
rect 240546 398898 240782 399134
rect 249546 399218 249782 399454
rect 249546 398898 249782 399134
rect 258546 399218 258782 399454
rect 258546 398898 258782 399134
rect 267546 399218 267782 399454
rect 267546 398898 267782 399134
rect 269348 399218 269584 399454
rect 269348 398898 269584 399134
rect 270720 399218 270956 399454
rect 270720 398898 270956 399134
rect 271566 399218 271802 399454
rect 271566 398898 271802 399134
rect 280566 399218 280802 399454
rect 280566 398898 280802 399134
rect 289566 399218 289802 399454
rect 289566 398898 289802 399134
rect 298566 399218 298802 399454
rect 298566 398898 298802 399134
rect 307566 399218 307802 399454
rect 307566 398898 307802 399134
rect 309368 399218 309604 399454
rect 309368 398898 309604 399134
rect 311740 399218 311976 399454
rect 311740 398898 311976 399134
rect 312586 399218 312822 399454
rect 312586 398898 312822 399134
rect 321586 399218 321822 399454
rect 321586 398898 321822 399134
rect 330586 399218 330822 399454
rect 330586 398898 330822 399134
rect 339586 399218 339822 399454
rect 339586 398898 339822 399134
rect 348586 399218 348822 399454
rect 348586 398898 348822 399134
rect 350388 399218 350624 399454
rect 350388 398898 350624 399134
rect 352760 399218 352996 399454
rect 352760 398898 352996 399134
rect 353606 399218 353842 399454
rect 353606 398898 353842 399134
rect 362606 399218 362842 399454
rect 362606 398898 362842 399134
rect 371606 399218 371842 399454
rect 371606 398898 371842 399134
rect 380606 399218 380842 399454
rect 380606 398898 380842 399134
rect 389606 399218 389842 399454
rect 389606 398898 389842 399134
rect 391408 399218 391644 399454
rect 391408 398898 391644 399134
rect 392780 399218 393016 399454
rect 392780 398898 393016 399134
rect 393626 399218 393862 399454
rect 393626 398898 393862 399134
rect 402626 399218 402862 399454
rect 402626 398898 402862 399134
rect 411626 399218 411862 399454
rect 411626 398898 411862 399134
rect 420626 399218 420862 399454
rect 420626 398898 420862 399134
rect 429626 399218 429862 399454
rect 429626 398898 429862 399134
rect 431428 399218 431664 399454
rect 431428 398898 431664 399134
rect 432800 399218 433036 399454
rect 432800 398898 433036 399134
rect 433646 399218 433882 399454
rect 433646 398898 433882 399134
rect 439432 399218 439668 399454
rect 439432 398898 439668 399134
rect 456610 399218 456846 399454
rect 456610 398898 456846 399134
rect 463442 399218 463678 399454
rect 463442 398898 463678 399134
rect 470648 399218 470884 399454
rect 470648 398898 470884 399134
rect 479648 399218 479884 399454
rect 479648 398898 479884 399134
rect 488648 399218 488884 399454
rect 488648 398898 488884 399134
rect 497648 399218 497884 399454
rect 497648 398898 497884 399134
rect 506648 399218 506884 399454
rect 506648 398898 506884 399134
rect 515648 399218 515884 399454
rect 515648 398898 515884 399134
rect 524648 399218 524884 399454
rect 524648 398898 524884 399134
rect 533648 399218 533884 399454
rect 533648 398898 533884 399134
rect 542648 399218 542884 399454
rect 542648 398898 542884 399134
rect 551648 399218 551884 399454
rect 551648 398898 551884 399134
rect 560648 399218 560884 399454
rect 560648 398898 560884 399134
rect 569648 399218 569884 399454
rect 569648 398898 569884 399134
rect 570850 399218 571086 399454
rect 570850 398898 571086 399134
rect 578670 399218 578906 399454
rect 578670 398898 578906 399134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 4582 381218 4818 381454
rect 4582 380898 4818 381134
rect 127058 381218 127294 381454
rect 127058 380898 127294 381134
rect 140296 381218 140532 381454
rect 140296 380898 140532 381134
rect 141102 381218 141338 381454
rect 141102 380898 141338 381134
rect 147648 381218 147884 381454
rect 147648 380898 147884 381134
rect 149300 381218 149536 381454
rect 149300 380898 149536 381134
rect 150106 381218 150342 381454
rect 150106 380898 150342 381134
rect 159106 381218 159342 381454
rect 159106 380898 159342 381134
rect 168106 381218 168342 381454
rect 168106 380898 168342 381134
rect 177106 381218 177342 381454
rect 177106 380898 177342 381134
rect 186106 381218 186342 381454
rect 186106 380898 186342 381134
rect 188668 381218 188904 381454
rect 188668 380898 188904 381134
rect 190320 381218 190556 381454
rect 190320 380898 190556 381134
rect 191126 381218 191362 381454
rect 191126 380898 191362 381134
rect 200126 381218 200362 381454
rect 200126 380898 200362 381134
rect 209126 381218 209362 381454
rect 209126 380898 209362 381134
rect 218126 381218 218362 381454
rect 218126 380898 218362 381134
rect 227126 381218 227362 381454
rect 227126 380898 227362 381134
rect 229688 381218 229924 381454
rect 229688 380898 229924 381134
rect 230340 381218 230576 381454
rect 230340 380898 230576 381134
rect 231146 381218 231382 381454
rect 231146 380898 231382 381134
rect 240146 381218 240382 381454
rect 240146 380898 240382 381134
rect 249146 381218 249382 381454
rect 249146 380898 249382 381134
rect 258146 381218 258382 381454
rect 258146 380898 258382 381134
rect 267146 381218 267382 381454
rect 267146 380898 267382 381134
rect 269708 381218 269944 381454
rect 269708 380898 269944 381134
rect 270360 381218 270596 381454
rect 270360 380898 270596 381134
rect 271166 381218 271402 381454
rect 271166 380898 271402 381134
rect 280166 381218 280402 381454
rect 280166 380898 280402 381134
rect 289166 381218 289402 381454
rect 289166 380898 289402 381134
rect 298166 381218 298402 381454
rect 298166 380898 298402 381134
rect 307166 381218 307402 381454
rect 307166 380898 307402 381134
rect 309728 381218 309964 381454
rect 309728 380898 309964 381134
rect 311380 381218 311616 381454
rect 311380 380898 311616 381134
rect 312186 381218 312422 381454
rect 312186 380898 312422 381134
rect 321186 381218 321422 381454
rect 321186 380898 321422 381134
rect 330186 381218 330422 381454
rect 330186 380898 330422 381134
rect 339186 381218 339422 381454
rect 339186 380898 339422 381134
rect 348186 381218 348422 381454
rect 348186 380898 348422 381134
rect 350748 381218 350984 381454
rect 350748 380898 350984 381134
rect 352400 381218 352636 381454
rect 352400 380898 352636 381134
rect 353206 381218 353442 381454
rect 353206 380898 353442 381134
rect 362206 381218 362442 381454
rect 362206 380898 362442 381134
rect 371206 381218 371442 381454
rect 371206 380898 371442 381134
rect 380206 381218 380442 381454
rect 380206 380898 380442 381134
rect 389206 381218 389442 381454
rect 389206 380898 389442 381134
rect 391768 381218 392004 381454
rect 391768 380898 392004 381134
rect 392420 381218 392656 381454
rect 392420 380898 392656 381134
rect 393226 381218 393462 381454
rect 393226 380898 393462 381134
rect 402226 381218 402462 381454
rect 402226 380898 402462 381134
rect 411226 381218 411462 381454
rect 411226 380898 411462 381134
rect 420226 381218 420462 381454
rect 420226 380898 420462 381134
rect 429226 381218 429462 381454
rect 429226 380898 429462 381134
rect 431788 381218 432024 381454
rect 431788 380898 432024 381134
rect 432440 381218 432676 381454
rect 432440 380898 432676 381134
rect 433246 381218 433482 381454
rect 433246 380898 433482 381134
rect 439792 381218 440028 381454
rect 439792 380898 440028 381134
rect 457010 381218 457246 381454
rect 457010 380898 457246 381134
rect 579470 381218 579706 381454
rect 579470 380898 579706 381134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect 5382 363218 5618 363454
rect 5382 362898 5618 363134
rect 127458 363218 127694 363454
rect 127458 362898 127694 363134
rect 140656 363218 140892 363454
rect 140656 362898 140892 363134
rect 141502 363218 141738 363454
rect 141502 362898 141738 363134
rect 147288 363218 147524 363454
rect 147288 362898 147524 363134
rect 149660 363218 149896 363454
rect 149660 362898 149896 363134
rect 150506 363218 150742 363454
rect 150506 362898 150742 363134
rect 159506 363218 159742 363454
rect 159506 362898 159742 363134
rect 168506 363218 168742 363454
rect 168506 362898 168742 363134
rect 177506 363218 177742 363454
rect 177506 362898 177742 363134
rect 186506 363218 186742 363454
rect 186506 362898 186742 363134
rect 188308 363218 188544 363454
rect 188308 362898 188544 363134
rect 190680 363218 190916 363454
rect 190680 362898 190916 363134
rect 191526 363218 191762 363454
rect 191526 362898 191762 363134
rect 200526 363218 200762 363454
rect 200526 362898 200762 363134
rect 209526 363218 209762 363454
rect 209526 362898 209762 363134
rect 218526 363218 218762 363454
rect 218526 362898 218762 363134
rect 227526 363218 227762 363454
rect 227526 362898 227762 363134
rect 229328 363218 229564 363454
rect 229328 362898 229564 363134
rect 230700 363218 230936 363454
rect 230700 362898 230936 363134
rect 231546 363218 231782 363454
rect 231546 362898 231782 363134
rect 240546 363218 240782 363454
rect 240546 362898 240782 363134
rect 249546 363218 249782 363454
rect 249546 362898 249782 363134
rect 258546 363218 258782 363454
rect 258546 362898 258782 363134
rect 267546 363218 267782 363454
rect 267546 362898 267782 363134
rect 269348 363218 269584 363454
rect 269348 362898 269584 363134
rect 270720 363218 270956 363454
rect 270720 362898 270956 363134
rect 271566 363218 271802 363454
rect 271566 362898 271802 363134
rect 280566 363218 280802 363454
rect 280566 362898 280802 363134
rect 289566 363218 289802 363454
rect 289566 362898 289802 363134
rect 298566 363218 298802 363454
rect 298566 362898 298802 363134
rect 307566 363218 307802 363454
rect 307566 362898 307802 363134
rect 309368 363218 309604 363454
rect 309368 362898 309604 363134
rect 311740 363218 311976 363454
rect 311740 362898 311976 363134
rect 312586 363218 312822 363454
rect 312586 362898 312822 363134
rect 321586 363218 321822 363454
rect 321586 362898 321822 363134
rect 330586 363218 330822 363454
rect 330586 362898 330822 363134
rect 339586 363218 339822 363454
rect 339586 362898 339822 363134
rect 348586 363218 348822 363454
rect 348586 362898 348822 363134
rect 350388 363218 350624 363454
rect 350388 362898 350624 363134
rect 352760 363218 352996 363454
rect 352760 362898 352996 363134
rect 353606 363218 353842 363454
rect 353606 362898 353842 363134
rect 362606 363218 362842 363454
rect 362606 362898 362842 363134
rect 371606 363218 371842 363454
rect 371606 362898 371842 363134
rect 380606 363218 380842 363454
rect 380606 362898 380842 363134
rect 389606 363218 389842 363454
rect 389606 362898 389842 363134
rect 391408 363218 391644 363454
rect 391408 362898 391644 363134
rect 392780 363218 393016 363454
rect 392780 362898 393016 363134
rect 393626 363218 393862 363454
rect 393626 362898 393862 363134
rect 402626 363218 402862 363454
rect 402626 362898 402862 363134
rect 411626 363218 411862 363454
rect 411626 362898 411862 363134
rect 420626 363218 420862 363454
rect 420626 362898 420862 363134
rect 429626 363218 429862 363454
rect 429626 362898 429862 363134
rect 431428 363218 431664 363454
rect 431428 362898 431664 363134
rect 432800 363218 433036 363454
rect 432800 362898 433036 363134
rect 433646 363218 433882 363454
rect 433646 362898 433882 363134
rect 439432 363218 439668 363454
rect 439432 362898 439668 363134
rect 456610 363218 456846 363454
rect 456610 362898 456846 363134
rect 578670 363218 578906 363454
rect 578670 362898 578906 363134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 4582 345218 4818 345454
rect 4582 344898 4818 345134
rect 127058 345218 127294 345454
rect 127058 344898 127294 345134
rect 140296 345218 140532 345454
rect 140296 344898 140532 345134
rect 141102 345218 141338 345454
rect 141102 344898 141338 345134
rect 147648 345218 147884 345454
rect 147648 344898 147884 345134
rect 149300 345218 149536 345454
rect 149300 344898 149536 345134
rect 150106 345218 150342 345454
rect 150106 344898 150342 345134
rect 159106 345218 159342 345454
rect 159106 344898 159342 345134
rect 168106 345218 168342 345454
rect 168106 344898 168342 345134
rect 177106 345218 177342 345454
rect 177106 344898 177342 345134
rect 186106 345218 186342 345454
rect 186106 344898 186342 345134
rect 188668 345218 188904 345454
rect 188668 344898 188904 345134
rect 190320 345218 190556 345454
rect 190320 344898 190556 345134
rect 191126 345218 191362 345454
rect 191126 344898 191362 345134
rect 200126 345218 200362 345454
rect 200126 344898 200362 345134
rect 209126 345218 209362 345454
rect 209126 344898 209362 345134
rect 218126 345218 218362 345454
rect 218126 344898 218362 345134
rect 227126 345218 227362 345454
rect 227126 344898 227362 345134
rect 229688 345218 229924 345454
rect 229688 344898 229924 345134
rect 230340 345218 230576 345454
rect 230340 344898 230576 345134
rect 231146 345218 231382 345454
rect 231146 344898 231382 345134
rect 240146 345218 240382 345454
rect 240146 344898 240382 345134
rect 249146 345218 249382 345454
rect 249146 344898 249382 345134
rect 258146 345218 258382 345454
rect 258146 344898 258382 345134
rect 267146 345218 267382 345454
rect 267146 344898 267382 345134
rect 269708 345218 269944 345454
rect 269708 344898 269944 345134
rect 270360 345218 270596 345454
rect 270360 344898 270596 345134
rect 271166 345218 271402 345454
rect 271166 344898 271402 345134
rect 280166 345218 280402 345454
rect 280166 344898 280402 345134
rect 289166 345218 289402 345454
rect 289166 344898 289402 345134
rect 298166 345218 298402 345454
rect 298166 344898 298402 345134
rect 307166 345218 307402 345454
rect 307166 344898 307402 345134
rect 309728 345218 309964 345454
rect 309728 344898 309964 345134
rect 311380 345218 311616 345454
rect 311380 344898 311616 345134
rect 312186 345218 312422 345454
rect 312186 344898 312422 345134
rect 321186 345218 321422 345454
rect 321186 344898 321422 345134
rect 330186 345218 330422 345454
rect 330186 344898 330422 345134
rect 339186 345218 339422 345454
rect 339186 344898 339422 345134
rect 348186 345218 348422 345454
rect 348186 344898 348422 345134
rect 350748 345218 350984 345454
rect 350748 344898 350984 345134
rect 352400 345218 352636 345454
rect 352400 344898 352636 345134
rect 353206 345218 353442 345454
rect 353206 344898 353442 345134
rect 362206 345218 362442 345454
rect 362206 344898 362442 345134
rect 371206 345218 371442 345454
rect 371206 344898 371442 345134
rect 380206 345218 380442 345454
rect 380206 344898 380442 345134
rect 389206 345218 389442 345454
rect 389206 344898 389442 345134
rect 391768 345218 392004 345454
rect 391768 344898 392004 345134
rect 392420 345218 392656 345454
rect 392420 344898 392656 345134
rect 393226 345218 393462 345454
rect 393226 344898 393462 345134
rect 402226 345218 402462 345454
rect 402226 344898 402462 345134
rect 411226 345218 411462 345454
rect 411226 344898 411462 345134
rect 420226 345218 420462 345454
rect 420226 344898 420462 345134
rect 429226 345218 429462 345454
rect 429226 344898 429462 345134
rect 431788 345218 432024 345454
rect 431788 344898 432024 345134
rect 432440 345218 432676 345454
rect 432440 344898 432676 345134
rect 433246 345218 433482 345454
rect 433246 344898 433482 345134
rect 439792 345218 440028 345454
rect 439792 344898 440028 345134
rect 457010 345218 457246 345454
rect 457010 344898 457246 345134
rect 579470 345218 579706 345454
rect 579470 344898 579706 345134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect 5382 327218 5618 327454
rect 5382 326898 5618 327134
rect 127458 327218 127694 327454
rect 127458 326898 127694 327134
rect 140656 327218 140892 327454
rect 140656 326898 140892 327134
rect 141502 327218 141738 327454
rect 141502 326898 141738 327134
rect 147288 327218 147524 327454
rect 147288 326898 147524 327134
rect 149660 327218 149896 327454
rect 149660 326898 149896 327134
rect 150506 327218 150742 327454
rect 150506 326898 150742 327134
rect 159506 327218 159742 327454
rect 159506 326898 159742 327134
rect 168506 327218 168742 327454
rect 168506 326898 168742 327134
rect 177506 327218 177742 327454
rect 177506 326898 177742 327134
rect 186506 327218 186742 327454
rect 186506 326898 186742 327134
rect 188308 327218 188544 327454
rect 188308 326898 188544 327134
rect 189768 327218 190004 327454
rect 189768 326898 190004 327134
rect 190680 327218 190916 327454
rect 190680 326898 190916 327134
rect 191526 327218 191762 327454
rect 191526 326898 191762 327134
rect 200526 327218 200762 327454
rect 200526 326898 200762 327134
rect 209526 327218 209762 327454
rect 209526 326898 209762 327134
rect 218526 327218 218762 327454
rect 218526 326898 218762 327134
rect 227526 327218 227762 327454
rect 227526 326898 227762 327134
rect 229328 327218 229564 327454
rect 229328 326898 229564 327134
rect 230700 327218 230936 327454
rect 230700 326898 230936 327134
rect 231546 327218 231782 327454
rect 231546 326898 231782 327134
rect 240546 327218 240782 327454
rect 240546 326898 240782 327134
rect 249546 327218 249782 327454
rect 249546 326898 249782 327134
rect 258546 327218 258782 327454
rect 258546 326898 258782 327134
rect 267546 327218 267782 327454
rect 267546 326898 267782 327134
rect 269348 327218 269584 327454
rect 269348 326898 269584 327134
rect 270720 327218 270956 327454
rect 270720 326898 270956 327134
rect 271566 327218 271802 327454
rect 271566 326898 271802 327134
rect 280566 327218 280802 327454
rect 280566 326898 280802 327134
rect 289566 327218 289802 327454
rect 289566 326898 289802 327134
rect 298566 327218 298802 327454
rect 298566 326898 298802 327134
rect 307566 327218 307802 327454
rect 307566 326898 307802 327134
rect 309368 327218 309604 327454
rect 309368 326898 309604 327134
rect 311740 327218 311976 327454
rect 311740 326898 311976 327134
rect 312586 327218 312822 327454
rect 312586 326898 312822 327134
rect 321586 327218 321822 327454
rect 321586 326898 321822 327134
rect 330586 327218 330822 327454
rect 330586 326898 330822 327134
rect 339586 327218 339822 327454
rect 339586 326898 339822 327134
rect 348586 327218 348822 327454
rect 348586 326898 348822 327134
rect 350388 327218 350624 327454
rect 350388 326898 350624 327134
rect 352760 327218 352996 327454
rect 352760 326898 352996 327134
rect 353606 327218 353842 327454
rect 353606 326898 353842 327134
rect 362606 327218 362842 327454
rect 362606 326898 362842 327134
rect 371606 327218 371842 327454
rect 371606 326898 371842 327134
rect 380606 327218 380842 327454
rect 380606 326898 380842 327134
rect 389606 327218 389842 327454
rect 389606 326898 389842 327134
rect 391408 327218 391644 327454
rect 391408 326898 391644 327134
rect 392780 327218 393016 327454
rect 392780 326898 393016 327134
rect 393626 327218 393862 327454
rect 393626 326898 393862 327134
rect 402626 327218 402862 327454
rect 402626 326898 402862 327134
rect 411626 327218 411862 327454
rect 411626 326898 411862 327134
rect 420626 327218 420862 327454
rect 420626 326898 420862 327134
rect 429626 327218 429862 327454
rect 429626 326898 429862 327134
rect 431428 327218 431664 327454
rect 431428 326898 431664 327134
rect 432800 327218 433036 327454
rect 432800 326898 433036 327134
rect 433646 327218 433882 327454
rect 433646 326898 433882 327134
rect 439432 327218 439668 327454
rect 439432 326898 439668 327134
rect 456610 327218 456846 327454
rect 456610 326898 456846 327134
rect 578670 327218 578906 327454
rect 578670 326898 578906 327134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 4582 309218 4818 309454
rect 4582 308898 4818 309134
rect 127058 309218 127294 309454
rect 127058 308898 127294 309134
rect 140296 309218 140532 309454
rect 140296 308898 140532 309134
rect 141102 309218 141338 309454
rect 141102 308898 141338 309134
rect 147648 309218 147884 309454
rect 147648 308898 147884 309134
rect 149300 309218 149536 309454
rect 149300 308898 149536 309134
rect 150106 309218 150342 309454
rect 150106 308898 150342 309134
rect 159106 309218 159342 309454
rect 159106 308898 159342 309134
rect 168106 309218 168342 309454
rect 168106 308898 168342 309134
rect 177106 309218 177342 309454
rect 177106 308898 177342 309134
rect 186106 309218 186342 309454
rect 186106 308898 186342 309134
rect 188668 309218 188904 309454
rect 188668 308898 188904 309134
rect 190320 309218 190556 309454
rect 190320 308898 190556 309134
rect 191126 309218 191362 309454
rect 191126 308898 191362 309134
rect 200126 309218 200362 309454
rect 200126 308898 200362 309134
rect 209126 309218 209362 309454
rect 209126 308898 209362 309134
rect 218126 309218 218362 309454
rect 218126 308898 218362 309134
rect 227126 309218 227362 309454
rect 227126 308898 227362 309134
rect 229688 309218 229924 309454
rect 229688 308898 229924 309134
rect 230340 309218 230576 309454
rect 230340 308898 230576 309134
rect 231146 309218 231382 309454
rect 231146 308898 231382 309134
rect 240146 309218 240382 309454
rect 240146 308898 240382 309134
rect 249146 309218 249382 309454
rect 249146 308898 249382 309134
rect 258146 309218 258382 309454
rect 258146 308898 258382 309134
rect 267146 309218 267382 309454
rect 267146 308898 267382 309134
rect 269708 309218 269944 309454
rect 269708 308898 269944 309134
rect 270360 309218 270596 309454
rect 270360 308898 270596 309134
rect 271166 309218 271402 309454
rect 271166 308898 271402 309134
rect 280166 309218 280402 309454
rect 280166 308898 280402 309134
rect 289166 309218 289402 309454
rect 289166 308898 289402 309134
rect 298166 309218 298402 309454
rect 298166 308898 298402 309134
rect 307166 309218 307402 309454
rect 307166 308898 307402 309134
rect 309728 309218 309964 309454
rect 309728 308898 309964 309134
rect 311380 309218 311616 309454
rect 311380 308898 311616 309134
rect 312186 309218 312422 309454
rect 312186 308898 312422 309134
rect 321186 309218 321422 309454
rect 321186 308898 321422 309134
rect 330186 309218 330422 309454
rect 330186 308898 330422 309134
rect 339186 309218 339422 309454
rect 339186 308898 339422 309134
rect 348186 309218 348422 309454
rect 348186 308898 348422 309134
rect 350748 309218 350984 309454
rect 350748 308898 350984 309134
rect 352400 309218 352636 309454
rect 352400 308898 352636 309134
rect 353206 309218 353442 309454
rect 353206 308898 353442 309134
rect 362206 309218 362442 309454
rect 362206 308898 362442 309134
rect 371206 309218 371442 309454
rect 371206 308898 371442 309134
rect 380206 309218 380442 309454
rect 380206 308898 380442 309134
rect 389206 309218 389442 309454
rect 389206 308898 389442 309134
rect 391768 309218 392004 309454
rect 391768 308898 392004 309134
rect 392420 309218 392656 309454
rect 392420 308898 392656 309134
rect 393226 309218 393462 309454
rect 393226 308898 393462 309134
rect 402226 309218 402462 309454
rect 402226 308898 402462 309134
rect 411226 309218 411462 309454
rect 411226 308898 411462 309134
rect 420226 309218 420462 309454
rect 420226 308898 420462 309134
rect 429226 309218 429462 309454
rect 429226 308898 429462 309134
rect 431788 309218 432024 309454
rect 431788 308898 432024 309134
rect 432440 309218 432676 309454
rect 432440 308898 432676 309134
rect 433246 309218 433482 309454
rect 433246 308898 433482 309134
rect 439792 309218 440028 309454
rect 439792 308898 440028 309134
rect 457010 309218 457246 309454
rect 457010 308898 457246 309134
rect 579470 309218 579706 309454
rect 579470 308898 579706 309134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect 5382 291218 5618 291454
rect 5382 290898 5618 291134
rect 108640 291218 108876 291454
rect 108640 290898 108876 291134
rect 109486 291218 109722 291454
rect 109486 290898 109722 291134
rect 118486 291218 118722 291454
rect 118486 290898 118722 291134
rect 127486 291218 127722 291454
rect 127486 290898 127722 291134
rect 136486 291218 136722 291454
rect 136486 290898 136722 291134
rect 145486 291218 145722 291454
rect 145486 290898 145722 291134
rect 147288 291218 147524 291454
rect 147288 290898 147524 291134
rect 149660 291218 149896 291454
rect 149660 290898 149896 291134
rect 150506 291218 150742 291454
rect 150506 290898 150742 291134
rect 159506 291218 159742 291454
rect 159506 290898 159742 291134
rect 168506 291218 168742 291454
rect 168506 290898 168742 291134
rect 177506 291218 177742 291454
rect 177506 290898 177742 291134
rect 186506 291218 186742 291454
rect 186506 290898 186742 291134
rect 188308 291218 188544 291454
rect 188308 290898 188544 291134
rect 190680 291218 190916 291454
rect 190680 290898 190916 291134
rect 191526 291218 191762 291454
rect 191526 290898 191762 291134
rect 200526 291218 200762 291454
rect 200526 290898 200762 291134
rect 209526 291218 209762 291454
rect 209526 290898 209762 291134
rect 218526 291218 218762 291454
rect 218526 290898 218762 291134
rect 227526 291218 227762 291454
rect 227526 290898 227762 291134
rect 229328 291218 229564 291454
rect 229328 290898 229564 291134
rect 230700 291218 230936 291454
rect 230700 290898 230936 291134
rect 231546 291218 231782 291454
rect 231546 290898 231782 291134
rect 240546 291218 240782 291454
rect 240546 290898 240782 291134
rect 249546 291218 249782 291454
rect 249546 290898 249782 291134
rect 258546 291218 258782 291454
rect 258546 290898 258782 291134
rect 267546 291218 267782 291454
rect 267546 290898 267782 291134
rect 269348 291218 269584 291454
rect 269348 290898 269584 291134
rect 270720 291218 270956 291454
rect 270720 290898 270956 291134
rect 271566 291218 271802 291454
rect 271566 290898 271802 291134
rect 280566 291218 280802 291454
rect 280566 290898 280802 291134
rect 289566 291218 289802 291454
rect 289566 290898 289802 291134
rect 298566 291218 298802 291454
rect 298566 290898 298802 291134
rect 307566 291218 307802 291454
rect 307566 290898 307802 291134
rect 309368 291218 309604 291454
rect 309368 290898 309604 291134
rect 311740 291218 311976 291454
rect 311740 290898 311976 291134
rect 312586 291218 312822 291454
rect 312586 290898 312822 291134
rect 321586 291218 321822 291454
rect 321586 290898 321822 291134
rect 330586 291218 330822 291454
rect 330586 290898 330822 291134
rect 339586 291218 339822 291454
rect 339586 290898 339822 291134
rect 348586 291218 348822 291454
rect 348586 290898 348822 291134
rect 350388 291218 350624 291454
rect 350388 290898 350624 291134
rect 352760 291218 352996 291454
rect 352760 290898 352996 291134
rect 353606 291218 353842 291454
rect 353606 290898 353842 291134
rect 362606 291218 362842 291454
rect 362606 290898 362842 291134
rect 371606 291218 371842 291454
rect 371606 290898 371842 291134
rect 380606 291218 380842 291454
rect 380606 290898 380842 291134
rect 389606 291218 389842 291454
rect 389606 290898 389842 291134
rect 391408 291218 391644 291454
rect 391408 290898 391644 291134
rect 392780 291218 393016 291454
rect 392780 290898 393016 291134
rect 393626 291218 393862 291454
rect 393626 290898 393862 291134
rect 402626 291218 402862 291454
rect 402626 290898 402862 291134
rect 411626 291218 411862 291454
rect 411626 290898 411862 291134
rect 420626 291218 420862 291454
rect 420626 290898 420862 291134
rect 429626 291218 429862 291454
rect 429626 290898 429862 291134
rect 431428 291218 431664 291454
rect 431428 290898 431664 291134
rect 432800 291218 433036 291454
rect 432800 290898 433036 291134
rect 433646 291218 433882 291454
rect 433646 290898 433882 291134
rect 442646 291218 442882 291454
rect 442646 290898 442882 291134
rect 451646 291218 451882 291454
rect 451646 290898 451882 291134
rect 460646 291218 460882 291454
rect 460646 290898 460882 291134
rect 469646 291218 469882 291454
rect 469646 290898 469882 291134
rect 471448 291218 471684 291454
rect 471448 290898 471684 291134
rect 578670 291218 578906 291454
rect 578670 290898 578906 291134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 4582 273218 4818 273454
rect 4582 272898 4818 273134
rect 108280 273218 108516 273454
rect 108280 272898 108516 273134
rect 109086 273218 109322 273454
rect 109086 272898 109322 273134
rect 118086 273218 118322 273454
rect 118086 272898 118322 273134
rect 127086 273218 127322 273454
rect 127086 272898 127322 273134
rect 136086 273218 136322 273454
rect 136086 272898 136322 273134
rect 145086 273218 145322 273454
rect 145086 272898 145322 273134
rect 147648 273218 147884 273454
rect 147648 272898 147884 273134
rect 148782 273218 149018 273454
rect 148782 272898 149018 273134
rect 149300 273218 149536 273454
rect 149300 272898 149536 273134
rect 150106 273218 150342 273454
rect 150106 272898 150342 273134
rect 159106 273218 159342 273454
rect 159106 272898 159342 273134
rect 168106 273218 168342 273454
rect 168106 272898 168342 273134
rect 177106 273218 177342 273454
rect 177106 272898 177342 273134
rect 186106 273218 186342 273454
rect 186106 272898 186342 273134
rect 188668 273218 188904 273454
rect 188668 272898 188904 273134
rect 189216 273218 189452 273454
rect 189216 272898 189452 273134
rect 190320 273218 190556 273454
rect 190320 272898 190556 273134
rect 191126 273218 191362 273454
rect 191126 272898 191362 273134
rect 200126 273218 200362 273454
rect 200126 272898 200362 273134
rect 209126 273218 209362 273454
rect 209126 272898 209362 273134
rect 218126 273218 218362 273454
rect 218126 272898 218362 273134
rect 227126 273218 227362 273454
rect 227126 272898 227362 273134
rect 229688 273218 229924 273454
rect 229688 272898 229924 273134
rect 230340 273218 230576 273454
rect 230340 272898 230576 273134
rect 231146 273218 231382 273454
rect 231146 272898 231382 273134
rect 240146 273218 240382 273454
rect 240146 272898 240382 273134
rect 249146 273218 249382 273454
rect 249146 272898 249382 273134
rect 258146 273218 258382 273454
rect 258146 272898 258382 273134
rect 267146 273218 267382 273454
rect 267146 272898 267382 273134
rect 269708 273218 269944 273454
rect 269708 272898 269944 273134
rect 270360 273218 270596 273454
rect 270360 272898 270596 273134
rect 271166 273218 271402 273454
rect 271166 272898 271402 273134
rect 280166 273218 280402 273454
rect 280166 272898 280402 273134
rect 289166 273218 289402 273454
rect 289166 272898 289402 273134
rect 298166 273218 298402 273454
rect 298166 272898 298402 273134
rect 307166 273218 307402 273454
rect 307166 272898 307402 273134
rect 309728 273218 309964 273454
rect 309728 272898 309964 273134
rect 310840 273218 311076 273454
rect 310840 272898 311076 273134
rect 311380 273218 311616 273454
rect 311380 272898 311616 273134
rect 312186 273218 312422 273454
rect 312186 272898 312422 273134
rect 321186 273218 321422 273454
rect 321186 272898 321422 273134
rect 330186 273218 330422 273454
rect 330186 272898 330422 273134
rect 339186 273218 339422 273454
rect 339186 272898 339422 273134
rect 348186 273218 348422 273454
rect 348186 272898 348422 273134
rect 350748 273218 350984 273454
rect 350748 272898 350984 273134
rect 351320 273218 351556 273454
rect 351320 272898 351556 273134
rect 352400 273218 352636 273454
rect 352400 272898 352636 273134
rect 353206 273218 353442 273454
rect 353206 272898 353442 273134
rect 362206 273218 362442 273454
rect 362206 272898 362442 273134
rect 371206 273218 371442 273454
rect 371206 272898 371442 273134
rect 380206 273218 380442 273454
rect 380206 272898 380442 273134
rect 389206 273218 389442 273454
rect 389206 272898 389442 273134
rect 391768 273218 392004 273454
rect 391768 272898 392004 273134
rect 392420 273218 392656 273454
rect 392420 272898 392656 273134
rect 393226 273218 393462 273454
rect 393226 272898 393462 273134
rect 402226 273218 402462 273454
rect 402226 272898 402462 273134
rect 411226 273218 411462 273454
rect 411226 272898 411462 273134
rect 420226 273218 420462 273454
rect 420226 272898 420462 273134
rect 429226 273218 429462 273454
rect 429226 272898 429462 273134
rect 431788 273218 432024 273454
rect 431788 272898 432024 273134
rect 432440 273218 432676 273454
rect 432440 272898 432676 273134
rect 433246 273218 433482 273454
rect 433246 272898 433482 273134
rect 442246 273218 442482 273454
rect 442246 272898 442482 273134
rect 451246 273218 451482 273454
rect 451246 272898 451482 273134
rect 460246 273218 460482 273454
rect 460246 272898 460482 273134
rect 469246 273218 469482 273454
rect 469246 272898 469482 273134
rect 471808 273218 472044 273454
rect 471808 272898 472044 273134
rect 579470 273218 579706 273454
rect 579470 272898 579706 273134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect 5382 255218 5618 255454
rect 5382 254898 5618 255134
rect 12592 255218 12828 255454
rect 12592 254898 12828 255134
rect 13438 255218 13674 255454
rect 13438 254898 13674 255134
rect 22438 255218 22674 255454
rect 22438 254898 22674 255134
rect 27228 255218 27464 255454
rect 27228 254898 27464 255134
rect 28600 255218 28836 255454
rect 28600 254898 28836 255134
rect 29446 255218 29682 255454
rect 29446 254898 29682 255134
rect 38446 255218 38682 255454
rect 38446 254898 38682 255134
rect 47446 255218 47682 255454
rect 47446 254898 47682 255134
rect 56446 255218 56682 255454
rect 56446 254898 56682 255134
rect 65446 255218 65682 255454
rect 65446 254898 65682 255134
rect 67248 255218 67484 255454
rect 67248 254898 67484 255134
rect 68620 255218 68856 255454
rect 68620 254898 68856 255134
rect 69466 255218 69702 255454
rect 69466 254898 69702 255134
rect 78466 255218 78702 255454
rect 78466 254898 78702 255134
rect 87466 255218 87702 255454
rect 87466 254898 87702 255134
rect 96466 255218 96702 255454
rect 96466 254898 96702 255134
rect 105466 255218 105702 255454
rect 105466 254898 105702 255134
rect 107268 255218 107504 255454
rect 107268 254898 107504 255134
rect 108640 255218 108876 255454
rect 108640 254898 108876 255134
rect 109486 255218 109722 255454
rect 109486 254898 109722 255134
rect 118486 255218 118722 255454
rect 118486 254898 118722 255134
rect 127486 255218 127722 255454
rect 127486 254898 127722 255134
rect 136486 255218 136722 255454
rect 136486 254898 136722 255134
rect 145486 255218 145722 255454
rect 145486 254898 145722 255134
rect 147288 255218 147524 255454
rect 147288 254898 147524 255134
rect 149660 255218 149896 255454
rect 149660 254898 149896 255134
rect 150506 255218 150742 255454
rect 150506 254898 150742 255134
rect 159506 255218 159742 255454
rect 159506 254898 159742 255134
rect 168506 255218 168742 255454
rect 168506 254898 168742 255134
rect 177506 255218 177742 255454
rect 177506 254898 177742 255134
rect 186506 255218 186742 255454
rect 186506 254898 186742 255134
rect 188308 255218 188544 255454
rect 188308 254898 188544 255134
rect 190680 255218 190916 255454
rect 190680 254898 190916 255134
rect 191526 255218 191762 255454
rect 191526 254898 191762 255134
rect 200526 255218 200762 255454
rect 200526 254898 200762 255134
rect 209526 255218 209762 255454
rect 209526 254898 209762 255134
rect 218526 255218 218762 255454
rect 218526 254898 218762 255134
rect 227526 255218 227762 255454
rect 227526 254898 227762 255134
rect 229328 255218 229564 255454
rect 229328 254898 229564 255134
rect 230700 255218 230936 255454
rect 230700 254898 230936 255134
rect 231546 255218 231782 255454
rect 231546 254898 231782 255134
rect 240546 255218 240782 255454
rect 240546 254898 240782 255134
rect 249546 255218 249782 255454
rect 249546 254898 249782 255134
rect 258546 255218 258782 255454
rect 258546 254898 258782 255134
rect 267546 255218 267782 255454
rect 267546 254898 267782 255134
rect 269348 255218 269584 255454
rect 269348 254898 269584 255134
rect 270720 255218 270956 255454
rect 270720 254898 270956 255134
rect 271566 255218 271802 255454
rect 271566 254898 271802 255134
rect 280566 255218 280802 255454
rect 280566 254898 280802 255134
rect 289566 255218 289802 255454
rect 289566 254898 289802 255134
rect 298566 255218 298802 255454
rect 298566 254898 298802 255134
rect 307566 255218 307802 255454
rect 307566 254898 307802 255134
rect 309368 255218 309604 255454
rect 309368 254898 309604 255134
rect 311740 255218 311976 255454
rect 311740 254898 311976 255134
rect 312586 255218 312822 255454
rect 312586 254898 312822 255134
rect 321586 255218 321822 255454
rect 321586 254898 321822 255134
rect 330586 255218 330822 255454
rect 330586 254898 330822 255134
rect 339586 255218 339822 255454
rect 339586 254898 339822 255134
rect 348586 255218 348822 255454
rect 348586 254898 348822 255134
rect 350388 255218 350624 255454
rect 350388 254898 350624 255134
rect 352760 255218 352996 255454
rect 352760 254898 352996 255134
rect 353606 255218 353842 255454
rect 353606 254898 353842 255134
rect 362606 255218 362842 255454
rect 362606 254898 362842 255134
rect 371606 255218 371842 255454
rect 371606 254898 371842 255134
rect 380606 255218 380842 255454
rect 380606 254898 380842 255134
rect 389606 255218 389842 255454
rect 389606 254898 389842 255134
rect 391408 255218 391644 255454
rect 391408 254898 391644 255134
rect 392780 255218 393016 255454
rect 392780 254898 393016 255134
rect 393626 255218 393862 255454
rect 393626 254898 393862 255134
rect 402626 255218 402862 255454
rect 402626 254898 402862 255134
rect 411626 255218 411862 255454
rect 411626 254898 411862 255134
rect 420626 255218 420862 255454
rect 420626 254898 420862 255134
rect 429626 255218 429862 255454
rect 429626 254898 429862 255134
rect 431428 255218 431664 255454
rect 431428 254898 431664 255134
rect 432800 255218 433036 255454
rect 432800 254898 433036 255134
rect 433646 255218 433882 255454
rect 433646 254898 433882 255134
rect 442646 255218 442882 255454
rect 442646 254898 442882 255134
rect 451646 255218 451882 255454
rect 451646 254898 451882 255134
rect 460646 255218 460882 255454
rect 460646 254898 460882 255134
rect 469646 255218 469882 255454
rect 469646 254898 469882 255134
rect 471448 255218 471684 255454
rect 471448 254898 471684 255134
rect 472820 255218 473056 255454
rect 472820 254898 473056 255134
rect 473666 255218 473902 255454
rect 473666 254898 473902 255134
rect 482666 255218 482902 255454
rect 482666 254898 482902 255134
rect 491666 255218 491902 255454
rect 491666 254898 491902 255134
rect 500666 255218 500902 255454
rect 500666 254898 500902 255134
rect 509666 255218 509902 255454
rect 509666 254898 509902 255134
rect 511468 255218 511704 255454
rect 511468 254898 511704 255134
rect 512840 255218 513076 255454
rect 512840 254898 513076 255134
rect 513686 255218 513922 255454
rect 513686 254898 513922 255134
rect 522686 255218 522922 255454
rect 522686 254898 522922 255134
rect 531686 255218 531922 255454
rect 531686 254898 531922 255134
rect 540686 255218 540922 255454
rect 540686 254898 540922 255134
rect 549686 255218 549922 255454
rect 549686 254898 549922 255134
rect 551488 255218 551724 255454
rect 551488 254898 551724 255134
rect 552860 255218 553096 255454
rect 552860 254898 553096 255134
rect 553706 255218 553942 255454
rect 553706 254898 553942 255134
rect 562706 255218 562942 255454
rect 562706 254898 562942 255134
rect 571706 255218 571942 255454
rect 571706 254898 571942 255134
rect 573476 255218 573712 255454
rect 573476 254898 573712 255134
rect 578670 255218 578906 255454
rect 578670 254898 578906 255134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 4582 237218 4818 237454
rect 4582 236898 4818 237134
rect 12232 237218 12468 237454
rect 12232 236898 12468 237134
rect 13038 237218 13274 237454
rect 13038 236898 13274 237134
rect 22038 237218 22274 237454
rect 22038 236898 22274 237134
rect 27588 237218 27824 237454
rect 27588 236898 27824 237134
rect 28240 237218 28476 237454
rect 28240 236898 28476 237134
rect 29046 237218 29282 237454
rect 29046 236898 29282 237134
rect 38046 237218 38282 237454
rect 38046 236898 38282 237134
rect 47046 237218 47282 237454
rect 47046 236898 47282 237134
rect 56046 237218 56282 237454
rect 56046 236898 56282 237134
rect 65046 237218 65282 237454
rect 65046 236898 65282 237134
rect 67608 237218 67844 237454
rect 67608 236898 67844 237134
rect 68260 237218 68496 237454
rect 68260 236898 68496 237134
rect 69066 237218 69302 237454
rect 69066 236898 69302 237134
rect 78066 237218 78302 237454
rect 78066 236898 78302 237134
rect 87066 237218 87302 237454
rect 87066 236898 87302 237134
rect 96066 237218 96302 237454
rect 96066 236898 96302 237134
rect 105066 237218 105302 237454
rect 105066 236898 105302 237134
rect 107628 237218 107864 237454
rect 107628 236898 107864 237134
rect 108280 237218 108516 237454
rect 108280 236898 108516 237134
rect 109086 237218 109322 237454
rect 109086 236898 109322 237134
rect 118086 237218 118322 237454
rect 118086 236898 118322 237134
rect 127086 237218 127322 237454
rect 127086 236898 127322 237134
rect 136086 237218 136322 237454
rect 136086 236898 136322 237134
rect 145086 237218 145322 237454
rect 145086 236898 145322 237134
rect 147648 237218 147884 237454
rect 147648 236898 147884 237134
rect 148782 237218 149018 237454
rect 148782 236898 149018 237134
rect 149300 237218 149536 237454
rect 149300 236898 149536 237134
rect 150106 237218 150342 237454
rect 150106 236898 150342 237134
rect 159106 237218 159342 237454
rect 159106 236898 159342 237134
rect 168106 237218 168342 237454
rect 168106 236898 168342 237134
rect 177106 237218 177342 237454
rect 177106 236898 177342 237134
rect 186106 237218 186342 237454
rect 186106 236898 186342 237134
rect 188668 237218 188904 237454
rect 188668 236898 188904 237134
rect 189216 237218 189452 237454
rect 189216 236898 189452 237134
rect 190320 237218 190556 237454
rect 190320 236898 190556 237134
rect 191126 237218 191362 237454
rect 191126 236898 191362 237134
rect 200126 237218 200362 237454
rect 200126 236898 200362 237134
rect 209126 237218 209362 237454
rect 209126 236898 209362 237134
rect 218126 237218 218362 237454
rect 218126 236898 218362 237134
rect 227126 237218 227362 237454
rect 227126 236898 227362 237134
rect 229688 237218 229924 237454
rect 229688 236898 229924 237134
rect 230340 237218 230576 237454
rect 230340 236898 230576 237134
rect 231146 237218 231382 237454
rect 231146 236898 231382 237134
rect 240146 237218 240382 237454
rect 240146 236898 240382 237134
rect 249146 237218 249382 237454
rect 249146 236898 249382 237134
rect 258146 237218 258382 237454
rect 258146 236898 258382 237134
rect 267146 237218 267382 237454
rect 267146 236898 267382 237134
rect 269708 237218 269944 237454
rect 269708 236898 269944 237134
rect 270360 237218 270596 237454
rect 270360 236898 270596 237134
rect 271166 237218 271402 237454
rect 271166 236898 271402 237134
rect 280166 237218 280402 237454
rect 280166 236898 280402 237134
rect 289166 237218 289402 237454
rect 289166 236898 289402 237134
rect 298166 237218 298402 237454
rect 298166 236898 298402 237134
rect 307166 237218 307402 237454
rect 307166 236898 307402 237134
rect 309728 237218 309964 237454
rect 309728 236898 309964 237134
rect 310840 237218 311076 237454
rect 310840 236898 311076 237134
rect 311380 237218 311616 237454
rect 311380 236898 311616 237134
rect 312186 237218 312422 237454
rect 312186 236898 312422 237134
rect 321186 237218 321422 237454
rect 321186 236898 321422 237134
rect 330186 237218 330422 237454
rect 330186 236898 330422 237134
rect 339186 237218 339422 237454
rect 339186 236898 339422 237134
rect 348186 237218 348422 237454
rect 348186 236898 348422 237134
rect 350748 237218 350984 237454
rect 350748 236898 350984 237134
rect 351320 237218 351556 237454
rect 351320 236898 351556 237134
rect 352400 237218 352636 237454
rect 352400 236898 352636 237134
rect 353206 237218 353442 237454
rect 353206 236898 353442 237134
rect 362206 237218 362442 237454
rect 362206 236898 362442 237134
rect 371206 237218 371442 237454
rect 371206 236898 371442 237134
rect 380206 237218 380442 237454
rect 380206 236898 380442 237134
rect 389206 237218 389442 237454
rect 389206 236898 389442 237134
rect 391768 237218 392004 237454
rect 391768 236898 392004 237134
rect 392420 237218 392656 237454
rect 392420 236898 392656 237134
rect 393226 237218 393462 237454
rect 393226 236898 393462 237134
rect 402226 237218 402462 237454
rect 402226 236898 402462 237134
rect 411226 237218 411462 237454
rect 411226 236898 411462 237134
rect 420226 237218 420462 237454
rect 420226 236898 420462 237134
rect 429226 237218 429462 237454
rect 429226 236898 429462 237134
rect 431788 237218 432024 237454
rect 431788 236898 432024 237134
rect 432440 237218 432676 237454
rect 432440 236898 432676 237134
rect 433246 237218 433482 237454
rect 433246 236898 433482 237134
rect 442246 237218 442482 237454
rect 442246 236898 442482 237134
rect 451246 237218 451482 237454
rect 451246 236898 451482 237134
rect 460246 237218 460482 237454
rect 460246 236898 460482 237134
rect 469246 237218 469482 237454
rect 469246 236898 469482 237134
rect 471808 237218 472044 237454
rect 471808 236898 472044 237134
rect 472460 237218 472696 237454
rect 472460 236898 472696 237134
rect 473266 237218 473502 237454
rect 473266 236898 473502 237134
rect 482266 237218 482502 237454
rect 482266 236898 482502 237134
rect 491266 237218 491502 237454
rect 491266 236898 491502 237134
rect 500266 237218 500502 237454
rect 500266 236898 500502 237134
rect 509266 237218 509502 237454
rect 509266 236898 509502 237134
rect 511828 237218 512064 237454
rect 511828 236898 512064 237134
rect 512480 237218 512716 237454
rect 512480 236898 512716 237134
rect 513286 237218 513522 237454
rect 513286 236898 513522 237134
rect 522286 237218 522522 237454
rect 522286 236898 522522 237134
rect 531286 237218 531522 237454
rect 531286 236898 531522 237134
rect 540286 237218 540522 237454
rect 540286 236898 540522 237134
rect 549286 237218 549522 237454
rect 549286 236898 549522 237134
rect 551848 237218 552084 237454
rect 551848 236898 552084 237134
rect 552500 237218 552736 237454
rect 552500 236898 552736 237134
rect 553306 237218 553542 237454
rect 553306 236898 553542 237134
rect 562306 237218 562542 237454
rect 562306 236898 562542 237134
rect 571306 237218 571542 237454
rect 571306 236898 571542 237134
rect 573836 237218 574072 237454
rect 573836 236898 574072 237134
rect 579470 237218 579706 237454
rect 579470 236898 579706 237134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect 5382 219218 5618 219454
rect 5382 218898 5618 219134
rect 12592 219218 12828 219454
rect 12592 218898 12828 219134
rect 13438 219218 13674 219454
rect 13438 218898 13674 219134
rect 22438 219218 22674 219454
rect 22438 218898 22674 219134
rect 27228 219218 27464 219454
rect 27228 218898 27464 219134
rect 28600 219218 28836 219454
rect 28600 218898 28836 219134
rect 29446 219218 29682 219454
rect 29446 218898 29682 219134
rect 38446 219218 38682 219454
rect 38446 218898 38682 219134
rect 47446 219218 47682 219454
rect 47446 218898 47682 219134
rect 56446 219218 56682 219454
rect 56446 218898 56682 219134
rect 65446 219218 65682 219454
rect 65446 218898 65682 219134
rect 67248 219218 67484 219454
rect 67248 218898 67484 219134
rect 68620 219218 68856 219454
rect 68620 218898 68856 219134
rect 69466 219218 69702 219454
rect 69466 218898 69702 219134
rect 78466 219218 78702 219454
rect 78466 218898 78702 219134
rect 87466 219218 87702 219454
rect 87466 218898 87702 219134
rect 96466 219218 96702 219454
rect 96466 218898 96702 219134
rect 105466 219218 105702 219454
rect 105466 218898 105702 219134
rect 107268 219218 107504 219454
rect 107268 218898 107504 219134
rect 108640 219218 108876 219454
rect 108640 218898 108876 219134
rect 109486 219218 109722 219454
rect 109486 218898 109722 219134
rect 118486 219218 118722 219454
rect 118486 218898 118722 219134
rect 127486 219218 127722 219454
rect 127486 218898 127722 219134
rect 136486 219218 136722 219454
rect 136486 218898 136722 219134
rect 145486 219218 145722 219454
rect 145486 218898 145722 219134
rect 147288 219218 147524 219454
rect 147288 218898 147524 219134
rect 149660 219218 149896 219454
rect 149660 218898 149896 219134
rect 150506 219218 150742 219454
rect 150506 218898 150742 219134
rect 159506 219218 159742 219454
rect 159506 218898 159742 219134
rect 168506 219218 168742 219454
rect 168506 218898 168742 219134
rect 177506 219218 177742 219454
rect 177506 218898 177742 219134
rect 186506 219218 186742 219454
rect 186506 218898 186742 219134
rect 188308 219218 188544 219454
rect 188308 218898 188544 219134
rect 190680 219218 190916 219454
rect 190680 218898 190916 219134
rect 191526 219218 191762 219454
rect 191526 218898 191762 219134
rect 200526 219218 200762 219454
rect 200526 218898 200762 219134
rect 209526 219218 209762 219454
rect 209526 218898 209762 219134
rect 218526 219218 218762 219454
rect 218526 218898 218762 219134
rect 227526 219218 227762 219454
rect 227526 218898 227762 219134
rect 229328 219218 229564 219454
rect 229328 218898 229564 219134
rect 230700 219218 230936 219454
rect 230700 218898 230936 219134
rect 231546 219218 231782 219454
rect 231546 218898 231782 219134
rect 240546 219218 240782 219454
rect 240546 218898 240782 219134
rect 249546 219218 249782 219454
rect 249546 218898 249782 219134
rect 258546 219218 258782 219454
rect 258546 218898 258782 219134
rect 267546 219218 267782 219454
rect 267546 218898 267782 219134
rect 269348 219218 269584 219454
rect 269348 218898 269584 219134
rect 270720 219218 270956 219454
rect 270720 218898 270956 219134
rect 271566 219218 271802 219454
rect 271566 218898 271802 219134
rect 280566 219218 280802 219454
rect 280566 218898 280802 219134
rect 289566 219218 289802 219454
rect 289566 218898 289802 219134
rect 298566 219218 298802 219454
rect 298566 218898 298802 219134
rect 307566 219218 307802 219454
rect 307566 218898 307802 219134
rect 309368 219218 309604 219454
rect 309368 218898 309604 219134
rect 311740 219218 311976 219454
rect 311740 218898 311976 219134
rect 312586 219218 312822 219454
rect 312586 218898 312822 219134
rect 321586 219218 321822 219454
rect 321586 218898 321822 219134
rect 330586 219218 330822 219454
rect 330586 218898 330822 219134
rect 339586 219218 339822 219454
rect 339586 218898 339822 219134
rect 348586 219218 348822 219454
rect 348586 218898 348822 219134
rect 350388 219218 350624 219454
rect 350388 218898 350624 219134
rect 352760 219218 352996 219454
rect 352760 218898 352996 219134
rect 353606 219218 353842 219454
rect 353606 218898 353842 219134
rect 362606 219218 362842 219454
rect 362606 218898 362842 219134
rect 371606 219218 371842 219454
rect 371606 218898 371842 219134
rect 380606 219218 380842 219454
rect 380606 218898 380842 219134
rect 389606 219218 389842 219454
rect 389606 218898 389842 219134
rect 391408 219218 391644 219454
rect 391408 218898 391644 219134
rect 392780 219218 393016 219454
rect 392780 218898 393016 219134
rect 393626 219218 393862 219454
rect 393626 218898 393862 219134
rect 402626 219218 402862 219454
rect 402626 218898 402862 219134
rect 411626 219218 411862 219454
rect 411626 218898 411862 219134
rect 420626 219218 420862 219454
rect 420626 218898 420862 219134
rect 429626 219218 429862 219454
rect 429626 218898 429862 219134
rect 431428 219218 431664 219454
rect 431428 218898 431664 219134
rect 432800 219218 433036 219454
rect 432800 218898 433036 219134
rect 433646 219218 433882 219454
rect 433646 218898 433882 219134
rect 442646 219218 442882 219454
rect 442646 218898 442882 219134
rect 451646 219218 451882 219454
rect 451646 218898 451882 219134
rect 460646 219218 460882 219454
rect 460646 218898 460882 219134
rect 469646 219218 469882 219454
rect 469646 218898 469882 219134
rect 471448 219218 471684 219454
rect 471448 218898 471684 219134
rect 472820 219218 473056 219454
rect 472820 218898 473056 219134
rect 473666 219218 473902 219454
rect 473666 218898 473902 219134
rect 482666 219218 482902 219454
rect 482666 218898 482902 219134
rect 491666 219218 491902 219454
rect 491666 218898 491902 219134
rect 500666 219218 500902 219454
rect 500666 218898 500902 219134
rect 509666 219218 509902 219454
rect 509666 218898 509902 219134
rect 511468 219218 511704 219454
rect 511468 218898 511704 219134
rect 512840 219218 513076 219454
rect 512840 218898 513076 219134
rect 513686 219218 513922 219454
rect 513686 218898 513922 219134
rect 522686 219218 522922 219454
rect 522686 218898 522922 219134
rect 531686 219218 531922 219454
rect 531686 218898 531922 219134
rect 540686 219218 540922 219454
rect 540686 218898 540922 219134
rect 549686 219218 549922 219454
rect 549686 218898 549922 219134
rect 551488 219218 551724 219454
rect 551488 218898 551724 219134
rect 552860 219218 553096 219454
rect 552860 218898 553096 219134
rect 553706 219218 553942 219454
rect 553706 218898 553942 219134
rect 562706 219218 562942 219454
rect 562706 218898 562942 219134
rect 571706 219218 571942 219454
rect 571706 218898 571942 219134
rect 573476 219218 573712 219454
rect 573476 218898 573712 219134
rect 578670 219218 578906 219454
rect 578670 218898 578906 219134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 4582 201218 4818 201454
rect 4582 200898 4818 201134
rect 12232 201218 12468 201454
rect 12232 200898 12468 201134
rect 13038 201218 13274 201454
rect 13038 200898 13274 201134
rect 22038 201218 22274 201454
rect 22038 200898 22274 201134
rect 27588 201218 27824 201454
rect 27588 200898 27824 201134
rect 28240 201218 28476 201454
rect 28240 200898 28476 201134
rect 29046 201218 29282 201454
rect 29046 200898 29282 201134
rect 38046 201218 38282 201454
rect 38046 200898 38282 201134
rect 47046 201218 47282 201454
rect 47046 200898 47282 201134
rect 56046 201218 56282 201454
rect 56046 200898 56282 201134
rect 65046 201218 65282 201454
rect 65046 200898 65282 201134
rect 67608 201218 67844 201454
rect 67608 200898 67844 201134
rect 68260 201218 68496 201454
rect 68260 200898 68496 201134
rect 69066 201218 69302 201454
rect 69066 200898 69302 201134
rect 78066 201218 78302 201454
rect 78066 200898 78302 201134
rect 87066 201218 87302 201454
rect 87066 200898 87302 201134
rect 96066 201218 96302 201454
rect 96066 200898 96302 201134
rect 105066 201218 105302 201454
rect 105066 200898 105302 201134
rect 107628 201218 107864 201454
rect 107628 200898 107864 201134
rect 108280 201218 108516 201454
rect 108280 200898 108516 201134
rect 109086 201218 109322 201454
rect 109086 200898 109322 201134
rect 118086 201218 118322 201454
rect 118086 200898 118322 201134
rect 127086 201218 127322 201454
rect 127086 200898 127322 201134
rect 136086 201218 136322 201454
rect 136086 200898 136322 201134
rect 145086 201218 145322 201454
rect 145086 200898 145322 201134
rect 147648 201218 147884 201454
rect 147648 200898 147884 201134
rect 149300 201218 149536 201454
rect 149300 200898 149536 201134
rect 150106 201218 150342 201454
rect 150106 200898 150342 201134
rect 159106 201218 159342 201454
rect 159106 200898 159342 201134
rect 168106 201218 168342 201454
rect 168106 200898 168342 201134
rect 177106 201218 177342 201454
rect 177106 200898 177342 201134
rect 186106 201218 186342 201454
rect 186106 200898 186342 201134
rect 188668 201218 188904 201454
rect 188668 200898 188904 201134
rect 190320 201218 190556 201454
rect 190320 200898 190556 201134
rect 191126 201218 191362 201454
rect 191126 200898 191362 201134
rect 200126 201218 200362 201454
rect 200126 200898 200362 201134
rect 209126 201218 209362 201454
rect 209126 200898 209362 201134
rect 218126 201218 218362 201454
rect 218126 200898 218362 201134
rect 227126 201218 227362 201454
rect 227126 200898 227362 201134
rect 229688 201218 229924 201454
rect 229688 200898 229924 201134
rect 230340 201218 230576 201454
rect 230340 200898 230576 201134
rect 231146 201218 231382 201454
rect 231146 200898 231382 201134
rect 240146 201218 240382 201454
rect 240146 200898 240382 201134
rect 249146 201218 249382 201454
rect 249146 200898 249382 201134
rect 258146 201218 258382 201454
rect 258146 200898 258382 201134
rect 267146 201218 267382 201454
rect 267146 200898 267382 201134
rect 269708 201218 269944 201454
rect 269708 200898 269944 201134
rect 270360 201218 270596 201454
rect 270360 200898 270596 201134
rect 271166 201218 271402 201454
rect 271166 200898 271402 201134
rect 280166 201218 280402 201454
rect 280166 200898 280402 201134
rect 289166 201218 289402 201454
rect 289166 200898 289402 201134
rect 298166 201218 298402 201454
rect 298166 200898 298402 201134
rect 307166 201218 307402 201454
rect 307166 200898 307402 201134
rect 309728 201218 309964 201454
rect 309728 200898 309964 201134
rect 311380 201218 311616 201454
rect 311380 200898 311616 201134
rect 312186 201218 312422 201454
rect 312186 200898 312422 201134
rect 321186 201218 321422 201454
rect 321186 200898 321422 201134
rect 330186 201218 330422 201454
rect 330186 200898 330422 201134
rect 339186 201218 339422 201454
rect 339186 200898 339422 201134
rect 348186 201218 348422 201454
rect 348186 200898 348422 201134
rect 350748 201218 350984 201454
rect 350748 200898 350984 201134
rect 352400 201218 352636 201454
rect 352400 200898 352636 201134
rect 353206 201218 353442 201454
rect 353206 200898 353442 201134
rect 362206 201218 362442 201454
rect 362206 200898 362442 201134
rect 371206 201218 371442 201454
rect 371206 200898 371442 201134
rect 380206 201218 380442 201454
rect 380206 200898 380442 201134
rect 389206 201218 389442 201454
rect 389206 200898 389442 201134
rect 391768 201218 392004 201454
rect 391768 200898 392004 201134
rect 392420 201218 392656 201454
rect 392420 200898 392656 201134
rect 393226 201218 393462 201454
rect 393226 200898 393462 201134
rect 402226 201218 402462 201454
rect 402226 200898 402462 201134
rect 411226 201218 411462 201454
rect 411226 200898 411462 201134
rect 420226 201218 420462 201454
rect 420226 200898 420462 201134
rect 429226 201218 429462 201454
rect 429226 200898 429462 201134
rect 431788 201218 432024 201454
rect 431788 200898 432024 201134
rect 432440 201218 432676 201454
rect 432440 200898 432676 201134
rect 433246 201218 433482 201454
rect 433246 200898 433482 201134
rect 442246 201218 442482 201454
rect 442246 200898 442482 201134
rect 451246 201218 451482 201454
rect 451246 200898 451482 201134
rect 460246 201218 460482 201454
rect 460246 200898 460482 201134
rect 469246 201218 469482 201454
rect 469246 200898 469482 201134
rect 471808 201218 472044 201454
rect 471808 200898 472044 201134
rect 472460 201218 472696 201454
rect 472460 200898 472696 201134
rect 473266 201218 473502 201454
rect 473266 200898 473502 201134
rect 482266 201218 482502 201454
rect 482266 200898 482502 201134
rect 491266 201218 491502 201454
rect 491266 200898 491502 201134
rect 500266 201218 500502 201454
rect 500266 200898 500502 201134
rect 509266 201218 509502 201454
rect 509266 200898 509502 201134
rect 511828 201218 512064 201454
rect 511828 200898 512064 201134
rect 512480 201218 512716 201454
rect 512480 200898 512716 201134
rect 513286 201218 513522 201454
rect 513286 200898 513522 201134
rect 522286 201218 522522 201454
rect 522286 200898 522522 201134
rect 531286 201218 531522 201454
rect 531286 200898 531522 201134
rect 540286 201218 540522 201454
rect 540286 200898 540522 201134
rect 549286 201218 549522 201454
rect 549286 200898 549522 201134
rect 551848 201218 552084 201454
rect 551848 200898 552084 201134
rect 552500 201218 552736 201454
rect 552500 200898 552736 201134
rect 553306 201218 553542 201454
rect 553306 200898 553542 201134
rect 562306 201218 562542 201454
rect 562306 200898 562542 201134
rect 571306 201218 571542 201454
rect 571306 200898 571542 201134
rect 573836 201218 574072 201454
rect 573836 200898 574072 201134
rect 579470 201218 579706 201454
rect 579470 200898 579706 201134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect 5382 183218 5618 183454
rect 5382 182898 5618 183134
rect 12592 183218 12828 183454
rect 12592 182898 12828 183134
rect 13438 183218 13674 183454
rect 13438 182898 13674 183134
rect 22438 183218 22674 183454
rect 22438 182898 22674 183134
rect 27228 183218 27464 183454
rect 27228 182898 27464 183134
rect 28600 183218 28836 183454
rect 28600 182898 28836 183134
rect 29446 183218 29682 183454
rect 29446 182898 29682 183134
rect 38446 183218 38682 183454
rect 38446 182898 38682 183134
rect 47446 183218 47682 183454
rect 47446 182898 47682 183134
rect 56446 183218 56682 183454
rect 56446 182898 56682 183134
rect 65446 183218 65682 183454
rect 65446 182898 65682 183134
rect 67248 183218 67484 183454
rect 67248 182898 67484 183134
rect 68620 183218 68856 183454
rect 68620 182898 68856 183134
rect 69466 183218 69702 183454
rect 69466 182898 69702 183134
rect 78466 183218 78702 183454
rect 78466 182898 78702 183134
rect 87466 183218 87702 183454
rect 87466 182898 87702 183134
rect 96466 183218 96702 183454
rect 96466 182898 96702 183134
rect 105466 183218 105702 183454
rect 105466 182898 105702 183134
rect 107268 183218 107504 183454
rect 107268 182898 107504 183134
rect 108640 183218 108876 183454
rect 108640 182898 108876 183134
rect 109486 183218 109722 183454
rect 109486 182898 109722 183134
rect 118486 183218 118722 183454
rect 118486 182898 118722 183134
rect 127486 183218 127722 183454
rect 127486 182898 127722 183134
rect 136486 183218 136722 183454
rect 136486 182898 136722 183134
rect 145486 183218 145722 183454
rect 145486 182898 145722 183134
rect 147288 183218 147524 183454
rect 147288 182898 147524 183134
rect 149660 183218 149896 183454
rect 149660 182898 149896 183134
rect 150506 183218 150742 183454
rect 150506 182898 150742 183134
rect 159506 183218 159742 183454
rect 159506 182898 159742 183134
rect 168506 183218 168742 183454
rect 168506 182898 168742 183134
rect 177506 183218 177742 183454
rect 177506 182898 177742 183134
rect 186506 183218 186742 183454
rect 186506 182898 186742 183134
rect 188308 183218 188544 183454
rect 188308 182898 188544 183134
rect 190680 183218 190916 183454
rect 190680 182898 190916 183134
rect 191526 183218 191762 183454
rect 191526 182898 191762 183134
rect 200526 183218 200762 183454
rect 200526 182898 200762 183134
rect 209526 183218 209762 183454
rect 209526 182898 209762 183134
rect 218526 183218 218762 183454
rect 218526 182898 218762 183134
rect 227526 183218 227762 183454
rect 227526 182898 227762 183134
rect 229328 183218 229564 183454
rect 229328 182898 229564 183134
rect 230700 183218 230936 183454
rect 230700 182898 230936 183134
rect 231546 183218 231782 183454
rect 231546 182898 231782 183134
rect 240546 183218 240782 183454
rect 240546 182898 240782 183134
rect 249546 183218 249782 183454
rect 249546 182898 249782 183134
rect 258546 183218 258782 183454
rect 258546 182898 258782 183134
rect 267546 183218 267782 183454
rect 267546 182898 267782 183134
rect 269348 183218 269584 183454
rect 269348 182898 269584 183134
rect 270720 183218 270956 183454
rect 270720 182898 270956 183134
rect 271566 183218 271802 183454
rect 271566 182898 271802 183134
rect 280566 183218 280802 183454
rect 280566 182898 280802 183134
rect 289566 183218 289802 183454
rect 289566 182898 289802 183134
rect 298566 183218 298802 183454
rect 298566 182898 298802 183134
rect 307566 183218 307802 183454
rect 307566 182898 307802 183134
rect 309368 183218 309604 183454
rect 309368 182898 309604 183134
rect 311740 183218 311976 183454
rect 311740 182898 311976 183134
rect 312586 183218 312822 183454
rect 312586 182898 312822 183134
rect 321586 183218 321822 183454
rect 321586 182898 321822 183134
rect 330586 183218 330822 183454
rect 330586 182898 330822 183134
rect 339586 183218 339822 183454
rect 339586 182898 339822 183134
rect 348586 183218 348822 183454
rect 348586 182898 348822 183134
rect 350388 183218 350624 183454
rect 350388 182898 350624 183134
rect 352760 183218 352996 183454
rect 352760 182898 352996 183134
rect 353606 183218 353842 183454
rect 353606 182898 353842 183134
rect 362606 183218 362842 183454
rect 362606 182898 362842 183134
rect 371606 183218 371842 183454
rect 371606 182898 371842 183134
rect 380606 183218 380842 183454
rect 380606 182898 380842 183134
rect 389606 183218 389842 183454
rect 389606 182898 389842 183134
rect 391408 183218 391644 183454
rect 391408 182898 391644 183134
rect 392780 183218 393016 183454
rect 392780 182898 393016 183134
rect 393626 183218 393862 183454
rect 393626 182898 393862 183134
rect 402626 183218 402862 183454
rect 402626 182898 402862 183134
rect 411626 183218 411862 183454
rect 411626 182898 411862 183134
rect 420626 183218 420862 183454
rect 420626 182898 420862 183134
rect 429626 183218 429862 183454
rect 429626 182898 429862 183134
rect 431428 183218 431664 183454
rect 431428 182898 431664 183134
rect 432800 183218 433036 183454
rect 432800 182898 433036 183134
rect 433646 183218 433882 183454
rect 433646 182898 433882 183134
rect 442646 183218 442882 183454
rect 442646 182898 442882 183134
rect 451646 183218 451882 183454
rect 451646 182898 451882 183134
rect 460646 183218 460882 183454
rect 460646 182898 460882 183134
rect 469646 183218 469882 183454
rect 469646 182898 469882 183134
rect 471448 183218 471684 183454
rect 471448 182898 471684 183134
rect 472820 183218 473056 183454
rect 472820 182898 473056 183134
rect 473666 183218 473902 183454
rect 473666 182898 473902 183134
rect 482666 183218 482902 183454
rect 482666 182898 482902 183134
rect 491666 183218 491902 183454
rect 491666 182898 491902 183134
rect 500666 183218 500902 183454
rect 500666 182898 500902 183134
rect 509666 183218 509902 183454
rect 509666 182898 509902 183134
rect 511468 183218 511704 183454
rect 511468 182898 511704 183134
rect 512840 183218 513076 183454
rect 512840 182898 513076 183134
rect 513686 183218 513922 183454
rect 513686 182898 513922 183134
rect 522686 183218 522922 183454
rect 522686 182898 522922 183134
rect 531686 183218 531922 183454
rect 531686 182898 531922 183134
rect 540686 183218 540922 183454
rect 540686 182898 540922 183134
rect 549686 183218 549922 183454
rect 549686 182898 549922 183134
rect 551488 183218 551724 183454
rect 551488 182898 551724 183134
rect 552860 183218 553096 183454
rect 552860 182898 553096 183134
rect 553706 183218 553942 183454
rect 553706 182898 553942 183134
rect 562706 183218 562942 183454
rect 562706 182898 562942 183134
rect 571706 183218 571942 183454
rect 571706 182898 571942 183134
rect 573476 183218 573712 183454
rect 573476 182898 573712 183134
rect 578670 183218 578906 183454
rect 578670 182898 578906 183134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 4582 165218 4818 165454
rect 4582 164898 4818 165134
rect 12232 165218 12468 165454
rect 12232 164898 12468 165134
rect 13038 165218 13274 165454
rect 13038 164898 13274 165134
rect 22038 165218 22274 165454
rect 22038 164898 22274 165134
rect 27588 165218 27824 165454
rect 27588 164898 27824 165134
rect 28240 165218 28476 165454
rect 28240 164898 28476 165134
rect 29046 165218 29282 165454
rect 29046 164898 29282 165134
rect 38046 165218 38282 165454
rect 38046 164898 38282 165134
rect 47046 165218 47282 165454
rect 47046 164898 47282 165134
rect 56046 165218 56282 165454
rect 56046 164898 56282 165134
rect 65046 165218 65282 165454
rect 65046 164898 65282 165134
rect 67608 165218 67844 165454
rect 67608 164898 67844 165134
rect 68260 165218 68496 165454
rect 68260 164898 68496 165134
rect 69066 165218 69302 165454
rect 69066 164898 69302 165134
rect 78066 165218 78302 165454
rect 78066 164898 78302 165134
rect 87066 165218 87302 165454
rect 87066 164898 87302 165134
rect 96066 165218 96302 165454
rect 96066 164898 96302 165134
rect 105066 165218 105302 165454
rect 105066 164898 105302 165134
rect 107628 165218 107864 165454
rect 107628 164898 107864 165134
rect 108280 165218 108516 165454
rect 108280 164898 108516 165134
rect 109086 165218 109322 165454
rect 109086 164898 109322 165134
rect 118086 165218 118322 165454
rect 118086 164898 118322 165134
rect 127086 165218 127322 165454
rect 127086 164898 127322 165134
rect 136086 165218 136322 165454
rect 136086 164898 136322 165134
rect 145086 165218 145322 165454
rect 145086 164898 145322 165134
rect 147648 165218 147884 165454
rect 147648 164898 147884 165134
rect 149300 165218 149536 165454
rect 149300 164898 149536 165134
rect 150106 165218 150342 165454
rect 150106 164898 150342 165134
rect 159106 165218 159342 165454
rect 159106 164898 159342 165134
rect 168106 165218 168342 165454
rect 168106 164898 168342 165134
rect 177106 165218 177342 165454
rect 177106 164898 177342 165134
rect 186106 165218 186342 165454
rect 186106 164898 186342 165134
rect 188668 165218 188904 165454
rect 188668 164898 188904 165134
rect 190320 165218 190556 165454
rect 190320 164898 190556 165134
rect 191126 165218 191362 165454
rect 191126 164898 191362 165134
rect 200126 165218 200362 165454
rect 200126 164898 200362 165134
rect 209126 165218 209362 165454
rect 209126 164898 209362 165134
rect 218126 165218 218362 165454
rect 218126 164898 218362 165134
rect 227126 165218 227362 165454
rect 227126 164898 227362 165134
rect 229688 165218 229924 165454
rect 229688 164898 229924 165134
rect 230340 165218 230576 165454
rect 230340 164898 230576 165134
rect 231146 165218 231382 165454
rect 231146 164898 231382 165134
rect 240146 165218 240382 165454
rect 240146 164898 240382 165134
rect 249146 165218 249382 165454
rect 249146 164898 249382 165134
rect 258146 165218 258382 165454
rect 258146 164898 258382 165134
rect 267146 165218 267382 165454
rect 267146 164898 267382 165134
rect 269708 165218 269944 165454
rect 269708 164898 269944 165134
rect 270360 165218 270596 165454
rect 270360 164898 270596 165134
rect 271166 165218 271402 165454
rect 271166 164898 271402 165134
rect 280166 165218 280402 165454
rect 280166 164898 280402 165134
rect 289166 165218 289402 165454
rect 289166 164898 289402 165134
rect 298166 165218 298402 165454
rect 298166 164898 298402 165134
rect 307166 165218 307402 165454
rect 307166 164898 307402 165134
rect 309728 165218 309964 165454
rect 309728 164898 309964 165134
rect 311380 165218 311616 165454
rect 311380 164898 311616 165134
rect 312186 165218 312422 165454
rect 312186 164898 312422 165134
rect 321186 165218 321422 165454
rect 321186 164898 321422 165134
rect 330186 165218 330422 165454
rect 330186 164898 330422 165134
rect 339186 165218 339422 165454
rect 339186 164898 339422 165134
rect 348186 165218 348422 165454
rect 348186 164898 348422 165134
rect 350748 165218 350984 165454
rect 350748 164898 350984 165134
rect 352400 165218 352636 165454
rect 352400 164898 352636 165134
rect 353206 165218 353442 165454
rect 353206 164898 353442 165134
rect 362206 165218 362442 165454
rect 362206 164898 362442 165134
rect 371206 165218 371442 165454
rect 371206 164898 371442 165134
rect 380206 165218 380442 165454
rect 380206 164898 380442 165134
rect 389206 165218 389442 165454
rect 389206 164898 389442 165134
rect 391768 165218 392004 165454
rect 391768 164898 392004 165134
rect 392420 165218 392656 165454
rect 392420 164898 392656 165134
rect 393226 165218 393462 165454
rect 393226 164898 393462 165134
rect 402226 165218 402462 165454
rect 402226 164898 402462 165134
rect 411226 165218 411462 165454
rect 411226 164898 411462 165134
rect 420226 165218 420462 165454
rect 420226 164898 420462 165134
rect 429226 165218 429462 165454
rect 429226 164898 429462 165134
rect 431788 165218 432024 165454
rect 431788 164898 432024 165134
rect 432440 165218 432676 165454
rect 432440 164898 432676 165134
rect 433246 165218 433482 165454
rect 433246 164898 433482 165134
rect 442246 165218 442482 165454
rect 442246 164898 442482 165134
rect 451246 165218 451482 165454
rect 451246 164898 451482 165134
rect 460246 165218 460482 165454
rect 460246 164898 460482 165134
rect 469246 165218 469482 165454
rect 469246 164898 469482 165134
rect 471808 165218 472044 165454
rect 471808 164898 472044 165134
rect 472460 165218 472696 165454
rect 472460 164898 472696 165134
rect 473266 165218 473502 165454
rect 473266 164898 473502 165134
rect 482266 165218 482502 165454
rect 482266 164898 482502 165134
rect 491266 165218 491502 165454
rect 491266 164898 491502 165134
rect 500266 165218 500502 165454
rect 500266 164898 500502 165134
rect 509266 165218 509502 165454
rect 509266 164898 509502 165134
rect 511828 165218 512064 165454
rect 511828 164898 512064 165134
rect 512480 165218 512716 165454
rect 512480 164898 512716 165134
rect 513286 165218 513522 165454
rect 513286 164898 513522 165134
rect 522286 165218 522522 165454
rect 522286 164898 522522 165134
rect 531286 165218 531522 165454
rect 531286 164898 531522 165134
rect 540286 165218 540522 165454
rect 540286 164898 540522 165134
rect 549286 165218 549522 165454
rect 549286 164898 549522 165134
rect 551848 165218 552084 165454
rect 551848 164898 552084 165134
rect 552500 165218 552736 165454
rect 552500 164898 552736 165134
rect 553306 165218 553542 165454
rect 553306 164898 553542 165134
rect 562306 165218 562542 165454
rect 562306 164898 562542 165134
rect 571306 165218 571542 165454
rect 571306 164898 571542 165134
rect 573836 165218 574072 165454
rect 573836 164898 574072 165134
rect 579470 165218 579706 165454
rect 579470 164898 579706 165134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect 5382 147218 5618 147454
rect 5382 146898 5618 147134
rect 12592 147218 12828 147454
rect 12592 146898 12828 147134
rect 13438 147218 13674 147454
rect 13438 146898 13674 147134
rect 22438 147218 22674 147454
rect 22438 146898 22674 147134
rect 27228 147218 27464 147454
rect 27228 146898 27464 147134
rect 28600 147218 28836 147454
rect 28600 146898 28836 147134
rect 29446 147218 29682 147454
rect 29446 146898 29682 147134
rect 38446 147218 38682 147454
rect 38446 146898 38682 147134
rect 47446 147218 47682 147454
rect 47446 146898 47682 147134
rect 56446 147218 56682 147454
rect 56446 146898 56682 147134
rect 65446 147218 65682 147454
rect 65446 146898 65682 147134
rect 67248 147218 67484 147454
rect 67248 146898 67484 147134
rect 68620 147218 68856 147454
rect 68620 146898 68856 147134
rect 69466 147218 69702 147454
rect 69466 146898 69702 147134
rect 78466 147218 78702 147454
rect 78466 146898 78702 147134
rect 87466 147218 87702 147454
rect 87466 146898 87702 147134
rect 96466 147218 96702 147454
rect 96466 146898 96702 147134
rect 105466 147218 105702 147454
rect 105466 146898 105702 147134
rect 107268 147218 107504 147454
rect 107268 146898 107504 147134
rect 108640 147218 108876 147454
rect 108640 146898 108876 147134
rect 109486 147218 109722 147454
rect 109486 146898 109722 147134
rect 118486 147218 118722 147454
rect 118486 146898 118722 147134
rect 127486 147218 127722 147454
rect 127486 146898 127722 147134
rect 136486 147218 136722 147454
rect 136486 146898 136722 147134
rect 145486 147218 145722 147454
rect 145486 146898 145722 147134
rect 147288 147218 147524 147454
rect 147288 146898 147524 147134
rect 149660 147218 149896 147454
rect 149660 146898 149896 147134
rect 150506 147218 150742 147454
rect 150506 146898 150742 147134
rect 159506 147218 159742 147454
rect 159506 146898 159742 147134
rect 168506 147218 168742 147454
rect 168506 146898 168742 147134
rect 177506 147218 177742 147454
rect 177506 146898 177742 147134
rect 186506 147218 186742 147454
rect 186506 146898 186742 147134
rect 188308 147218 188544 147454
rect 188308 146898 188544 147134
rect 190680 147218 190916 147454
rect 190680 146898 190916 147134
rect 191526 147218 191762 147454
rect 191526 146898 191762 147134
rect 200526 147218 200762 147454
rect 200526 146898 200762 147134
rect 209526 147218 209762 147454
rect 209526 146898 209762 147134
rect 218526 147218 218762 147454
rect 218526 146898 218762 147134
rect 227526 147218 227762 147454
rect 227526 146898 227762 147134
rect 229328 147218 229564 147454
rect 229328 146898 229564 147134
rect 230700 147218 230936 147454
rect 230700 146898 230936 147134
rect 231546 147218 231782 147454
rect 231546 146898 231782 147134
rect 240546 147218 240782 147454
rect 240546 146898 240782 147134
rect 249546 147218 249782 147454
rect 249546 146898 249782 147134
rect 258546 147218 258782 147454
rect 258546 146898 258782 147134
rect 267546 147218 267782 147454
rect 267546 146898 267782 147134
rect 269348 147218 269584 147454
rect 269348 146898 269584 147134
rect 270720 147218 270956 147454
rect 270720 146898 270956 147134
rect 271566 147218 271802 147454
rect 271566 146898 271802 147134
rect 280566 147218 280802 147454
rect 280566 146898 280802 147134
rect 289566 147218 289802 147454
rect 289566 146898 289802 147134
rect 298566 147218 298802 147454
rect 298566 146898 298802 147134
rect 307566 147218 307802 147454
rect 307566 146898 307802 147134
rect 309368 147218 309604 147454
rect 309368 146898 309604 147134
rect 311740 147218 311976 147454
rect 311740 146898 311976 147134
rect 312586 147218 312822 147454
rect 312586 146898 312822 147134
rect 321586 147218 321822 147454
rect 321586 146898 321822 147134
rect 330586 147218 330822 147454
rect 330586 146898 330822 147134
rect 339586 147218 339822 147454
rect 339586 146898 339822 147134
rect 348586 147218 348822 147454
rect 348586 146898 348822 147134
rect 350388 147218 350624 147454
rect 350388 146898 350624 147134
rect 352760 147218 352996 147454
rect 352760 146898 352996 147134
rect 353606 147218 353842 147454
rect 353606 146898 353842 147134
rect 362606 147218 362842 147454
rect 362606 146898 362842 147134
rect 371606 147218 371842 147454
rect 371606 146898 371842 147134
rect 380606 147218 380842 147454
rect 380606 146898 380842 147134
rect 389606 147218 389842 147454
rect 389606 146898 389842 147134
rect 391408 147218 391644 147454
rect 391408 146898 391644 147134
rect 392780 147218 393016 147454
rect 392780 146898 393016 147134
rect 393626 147218 393862 147454
rect 393626 146898 393862 147134
rect 402626 147218 402862 147454
rect 402626 146898 402862 147134
rect 411626 147218 411862 147454
rect 411626 146898 411862 147134
rect 420626 147218 420862 147454
rect 420626 146898 420862 147134
rect 429626 147218 429862 147454
rect 429626 146898 429862 147134
rect 431428 147218 431664 147454
rect 431428 146898 431664 147134
rect 432800 147218 433036 147454
rect 432800 146898 433036 147134
rect 433646 147218 433882 147454
rect 433646 146898 433882 147134
rect 442646 147218 442882 147454
rect 442646 146898 442882 147134
rect 451646 147218 451882 147454
rect 451646 146898 451882 147134
rect 460646 147218 460882 147454
rect 460646 146898 460882 147134
rect 469646 147218 469882 147454
rect 469646 146898 469882 147134
rect 471448 147218 471684 147454
rect 471448 146898 471684 147134
rect 472820 147218 473056 147454
rect 472820 146898 473056 147134
rect 473666 147218 473902 147454
rect 473666 146898 473902 147134
rect 482666 147218 482902 147454
rect 482666 146898 482902 147134
rect 491666 147218 491902 147454
rect 491666 146898 491902 147134
rect 500666 147218 500902 147454
rect 500666 146898 500902 147134
rect 509666 147218 509902 147454
rect 509666 146898 509902 147134
rect 511468 147218 511704 147454
rect 511468 146898 511704 147134
rect 512840 147218 513076 147454
rect 512840 146898 513076 147134
rect 513686 147218 513922 147454
rect 513686 146898 513922 147134
rect 522686 147218 522922 147454
rect 522686 146898 522922 147134
rect 531686 147218 531922 147454
rect 531686 146898 531922 147134
rect 540686 147218 540922 147454
rect 540686 146898 540922 147134
rect 549686 147218 549922 147454
rect 549686 146898 549922 147134
rect 551488 147218 551724 147454
rect 551488 146898 551724 147134
rect 552860 147218 553096 147454
rect 552860 146898 553096 147134
rect 553706 147218 553942 147454
rect 553706 146898 553942 147134
rect 562706 147218 562942 147454
rect 562706 146898 562942 147134
rect 571706 147218 571942 147454
rect 571706 146898 571942 147134
rect 573476 147218 573712 147454
rect 573476 146898 573712 147134
rect 578670 147218 578906 147454
rect 578670 146898 578906 147134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 4582 129218 4818 129454
rect 4582 128898 4818 129134
rect 12232 129218 12468 129454
rect 12232 128898 12468 129134
rect 13038 129218 13274 129454
rect 13038 128898 13274 129134
rect 22038 129218 22274 129454
rect 22038 128898 22274 129134
rect 27588 129218 27824 129454
rect 27588 128898 27824 129134
rect 28240 129218 28476 129454
rect 28240 128898 28476 129134
rect 29046 129218 29282 129454
rect 29046 128898 29282 129134
rect 38046 129218 38282 129454
rect 38046 128898 38282 129134
rect 47046 129218 47282 129454
rect 47046 128898 47282 129134
rect 56046 129218 56282 129454
rect 56046 128898 56282 129134
rect 65046 129218 65282 129454
rect 65046 128898 65282 129134
rect 67608 129218 67844 129454
rect 67608 128898 67844 129134
rect 68260 129218 68496 129454
rect 68260 128898 68496 129134
rect 69066 129218 69302 129454
rect 69066 128898 69302 129134
rect 78066 129218 78302 129454
rect 78066 128898 78302 129134
rect 87066 129218 87302 129454
rect 87066 128898 87302 129134
rect 96066 129218 96302 129454
rect 96066 128898 96302 129134
rect 105066 129218 105302 129454
rect 105066 128898 105302 129134
rect 107628 129218 107864 129454
rect 107628 128898 107864 129134
rect 108280 129218 108516 129454
rect 108280 128898 108516 129134
rect 109086 129218 109322 129454
rect 109086 128898 109322 129134
rect 118086 129218 118322 129454
rect 118086 128898 118322 129134
rect 127086 129218 127322 129454
rect 127086 128898 127322 129134
rect 136086 129218 136322 129454
rect 136086 128898 136322 129134
rect 145086 129218 145322 129454
rect 145086 128898 145322 129134
rect 147648 129218 147884 129454
rect 147648 128898 147884 129134
rect 149300 129218 149536 129454
rect 149300 128898 149536 129134
rect 150106 129218 150342 129454
rect 150106 128898 150342 129134
rect 159106 129218 159342 129454
rect 159106 128898 159342 129134
rect 168106 129218 168342 129454
rect 168106 128898 168342 129134
rect 177106 129218 177342 129454
rect 177106 128898 177342 129134
rect 186106 129218 186342 129454
rect 186106 128898 186342 129134
rect 188668 129218 188904 129454
rect 188668 128898 188904 129134
rect 190320 129218 190556 129454
rect 190320 128898 190556 129134
rect 191126 129218 191362 129454
rect 191126 128898 191362 129134
rect 200126 129218 200362 129454
rect 200126 128898 200362 129134
rect 209126 129218 209362 129454
rect 209126 128898 209362 129134
rect 218126 129218 218362 129454
rect 218126 128898 218362 129134
rect 227126 129218 227362 129454
rect 227126 128898 227362 129134
rect 229688 129218 229924 129454
rect 229688 128898 229924 129134
rect 230340 129218 230576 129454
rect 230340 128898 230576 129134
rect 231146 129218 231382 129454
rect 231146 128898 231382 129134
rect 240146 129218 240382 129454
rect 240146 128898 240382 129134
rect 249146 129218 249382 129454
rect 249146 128898 249382 129134
rect 258146 129218 258382 129454
rect 258146 128898 258382 129134
rect 267146 129218 267382 129454
rect 267146 128898 267382 129134
rect 269708 129218 269944 129454
rect 269708 128898 269944 129134
rect 270360 129218 270596 129454
rect 270360 128898 270596 129134
rect 271166 129218 271402 129454
rect 271166 128898 271402 129134
rect 280166 129218 280402 129454
rect 280166 128898 280402 129134
rect 289166 129218 289402 129454
rect 289166 128898 289402 129134
rect 298166 129218 298402 129454
rect 298166 128898 298402 129134
rect 307166 129218 307402 129454
rect 307166 128898 307402 129134
rect 309728 129218 309964 129454
rect 309728 128898 309964 129134
rect 311380 129218 311616 129454
rect 311380 128898 311616 129134
rect 312186 129218 312422 129454
rect 312186 128898 312422 129134
rect 321186 129218 321422 129454
rect 321186 128898 321422 129134
rect 330186 129218 330422 129454
rect 330186 128898 330422 129134
rect 339186 129218 339422 129454
rect 339186 128898 339422 129134
rect 348186 129218 348422 129454
rect 348186 128898 348422 129134
rect 350748 129218 350984 129454
rect 350748 128898 350984 129134
rect 352400 129218 352636 129454
rect 352400 128898 352636 129134
rect 353206 129218 353442 129454
rect 353206 128898 353442 129134
rect 362206 129218 362442 129454
rect 362206 128898 362442 129134
rect 371206 129218 371442 129454
rect 371206 128898 371442 129134
rect 380206 129218 380442 129454
rect 380206 128898 380442 129134
rect 389206 129218 389442 129454
rect 389206 128898 389442 129134
rect 391768 129218 392004 129454
rect 391768 128898 392004 129134
rect 392420 129218 392656 129454
rect 392420 128898 392656 129134
rect 393226 129218 393462 129454
rect 393226 128898 393462 129134
rect 402226 129218 402462 129454
rect 402226 128898 402462 129134
rect 411226 129218 411462 129454
rect 411226 128898 411462 129134
rect 420226 129218 420462 129454
rect 420226 128898 420462 129134
rect 429226 129218 429462 129454
rect 429226 128898 429462 129134
rect 431788 129218 432024 129454
rect 431788 128898 432024 129134
rect 432440 129218 432676 129454
rect 432440 128898 432676 129134
rect 433246 129218 433482 129454
rect 433246 128898 433482 129134
rect 442246 129218 442482 129454
rect 442246 128898 442482 129134
rect 451246 129218 451482 129454
rect 451246 128898 451482 129134
rect 460246 129218 460482 129454
rect 460246 128898 460482 129134
rect 469246 129218 469482 129454
rect 469246 128898 469482 129134
rect 471808 129218 472044 129454
rect 471808 128898 472044 129134
rect 472460 129218 472696 129454
rect 472460 128898 472696 129134
rect 473266 129218 473502 129454
rect 473266 128898 473502 129134
rect 482266 129218 482502 129454
rect 482266 128898 482502 129134
rect 491266 129218 491502 129454
rect 491266 128898 491502 129134
rect 500266 129218 500502 129454
rect 500266 128898 500502 129134
rect 509266 129218 509502 129454
rect 509266 128898 509502 129134
rect 511828 129218 512064 129454
rect 511828 128898 512064 129134
rect 512480 129218 512716 129454
rect 512480 128898 512716 129134
rect 513286 129218 513522 129454
rect 513286 128898 513522 129134
rect 522286 129218 522522 129454
rect 522286 128898 522522 129134
rect 531286 129218 531522 129454
rect 531286 128898 531522 129134
rect 540286 129218 540522 129454
rect 540286 128898 540522 129134
rect 549286 129218 549522 129454
rect 549286 128898 549522 129134
rect 551848 129218 552084 129454
rect 551848 128898 552084 129134
rect 552500 129218 552736 129454
rect 552500 128898 552736 129134
rect 553306 129218 553542 129454
rect 553306 128898 553542 129134
rect 562306 129218 562542 129454
rect 562306 128898 562542 129134
rect 571306 129218 571542 129454
rect 571306 128898 571542 129134
rect 573836 129218 574072 129454
rect 573836 128898 574072 129134
rect 579470 129218 579706 129454
rect 579470 128898 579706 129134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect 5382 111218 5618 111454
rect 5382 110898 5618 111134
rect 12592 111218 12828 111454
rect 12592 110898 12828 111134
rect 13438 111218 13674 111454
rect 13438 110898 13674 111134
rect 22438 111218 22674 111454
rect 22438 110898 22674 111134
rect 27228 111218 27464 111454
rect 27228 110898 27464 111134
rect 28600 111218 28836 111454
rect 28600 110898 28836 111134
rect 29446 111218 29682 111454
rect 29446 110898 29682 111134
rect 38446 111218 38682 111454
rect 38446 110898 38682 111134
rect 47446 111218 47682 111454
rect 47446 110898 47682 111134
rect 56446 111218 56682 111454
rect 56446 110898 56682 111134
rect 65446 111218 65682 111454
rect 65446 110898 65682 111134
rect 67248 111218 67484 111454
rect 67248 110898 67484 111134
rect 68620 111218 68856 111454
rect 68620 110898 68856 111134
rect 69466 111218 69702 111454
rect 69466 110898 69702 111134
rect 78466 111218 78702 111454
rect 78466 110898 78702 111134
rect 87466 111218 87702 111454
rect 87466 110898 87702 111134
rect 96466 111218 96702 111454
rect 96466 110898 96702 111134
rect 105466 111218 105702 111454
rect 105466 110898 105702 111134
rect 107268 111218 107504 111454
rect 107268 110898 107504 111134
rect 108640 111218 108876 111454
rect 108640 110898 108876 111134
rect 109486 111218 109722 111454
rect 109486 110898 109722 111134
rect 118486 111218 118722 111454
rect 118486 110898 118722 111134
rect 127486 111218 127722 111454
rect 127486 110898 127722 111134
rect 136486 111218 136722 111454
rect 136486 110898 136722 111134
rect 145486 111218 145722 111454
rect 145486 110898 145722 111134
rect 147288 111218 147524 111454
rect 147288 110898 147524 111134
rect 149660 111218 149896 111454
rect 149660 110898 149896 111134
rect 150506 111218 150742 111454
rect 150506 110898 150742 111134
rect 159506 111218 159742 111454
rect 159506 110898 159742 111134
rect 168506 111218 168742 111454
rect 168506 110898 168742 111134
rect 177506 111218 177742 111454
rect 177506 110898 177742 111134
rect 186506 111218 186742 111454
rect 186506 110898 186742 111134
rect 188308 111218 188544 111454
rect 188308 110898 188544 111134
rect 190680 111218 190916 111454
rect 190680 110898 190916 111134
rect 191526 111218 191762 111454
rect 191526 110898 191762 111134
rect 200526 111218 200762 111454
rect 200526 110898 200762 111134
rect 209526 111218 209762 111454
rect 209526 110898 209762 111134
rect 218526 111218 218762 111454
rect 218526 110898 218762 111134
rect 227526 111218 227762 111454
rect 227526 110898 227762 111134
rect 229328 111218 229564 111454
rect 229328 110898 229564 111134
rect 230700 111218 230936 111454
rect 230700 110898 230936 111134
rect 231546 111218 231782 111454
rect 231546 110898 231782 111134
rect 240546 111218 240782 111454
rect 240546 110898 240782 111134
rect 249546 111218 249782 111454
rect 249546 110898 249782 111134
rect 258546 111218 258782 111454
rect 258546 110898 258782 111134
rect 267546 111218 267782 111454
rect 267546 110898 267782 111134
rect 269348 111218 269584 111454
rect 269348 110898 269584 111134
rect 270720 111218 270956 111454
rect 270720 110898 270956 111134
rect 271566 111218 271802 111454
rect 271566 110898 271802 111134
rect 280566 111218 280802 111454
rect 280566 110898 280802 111134
rect 289566 111218 289802 111454
rect 289566 110898 289802 111134
rect 298566 111218 298802 111454
rect 298566 110898 298802 111134
rect 307566 111218 307802 111454
rect 307566 110898 307802 111134
rect 309368 111218 309604 111454
rect 309368 110898 309604 111134
rect 311740 111218 311976 111454
rect 311740 110898 311976 111134
rect 312586 111218 312822 111454
rect 312586 110898 312822 111134
rect 321586 111218 321822 111454
rect 321586 110898 321822 111134
rect 330586 111218 330822 111454
rect 330586 110898 330822 111134
rect 339586 111218 339822 111454
rect 339586 110898 339822 111134
rect 348586 111218 348822 111454
rect 348586 110898 348822 111134
rect 350388 111218 350624 111454
rect 350388 110898 350624 111134
rect 352760 111218 352996 111454
rect 352760 110898 352996 111134
rect 353606 111218 353842 111454
rect 353606 110898 353842 111134
rect 362606 111218 362842 111454
rect 362606 110898 362842 111134
rect 371606 111218 371842 111454
rect 371606 110898 371842 111134
rect 380606 111218 380842 111454
rect 380606 110898 380842 111134
rect 389606 111218 389842 111454
rect 389606 110898 389842 111134
rect 391408 111218 391644 111454
rect 391408 110898 391644 111134
rect 392780 111218 393016 111454
rect 392780 110898 393016 111134
rect 393626 111218 393862 111454
rect 393626 110898 393862 111134
rect 402626 111218 402862 111454
rect 402626 110898 402862 111134
rect 411626 111218 411862 111454
rect 411626 110898 411862 111134
rect 420626 111218 420862 111454
rect 420626 110898 420862 111134
rect 429626 111218 429862 111454
rect 429626 110898 429862 111134
rect 431428 111218 431664 111454
rect 431428 110898 431664 111134
rect 432800 111218 433036 111454
rect 432800 110898 433036 111134
rect 433646 111218 433882 111454
rect 433646 110898 433882 111134
rect 442646 111218 442882 111454
rect 442646 110898 442882 111134
rect 451646 111218 451882 111454
rect 451646 110898 451882 111134
rect 460646 111218 460882 111454
rect 460646 110898 460882 111134
rect 469646 111218 469882 111454
rect 469646 110898 469882 111134
rect 471448 111218 471684 111454
rect 471448 110898 471684 111134
rect 472820 111218 473056 111454
rect 472820 110898 473056 111134
rect 473666 111218 473902 111454
rect 473666 110898 473902 111134
rect 482666 111218 482902 111454
rect 482666 110898 482902 111134
rect 491666 111218 491902 111454
rect 491666 110898 491902 111134
rect 500666 111218 500902 111454
rect 500666 110898 500902 111134
rect 509666 111218 509902 111454
rect 509666 110898 509902 111134
rect 511468 111218 511704 111454
rect 511468 110898 511704 111134
rect 512840 111218 513076 111454
rect 512840 110898 513076 111134
rect 513686 111218 513922 111454
rect 513686 110898 513922 111134
rect 522686 111218 522922 111454
rect 522686 110898 522922 111134
rect 531686 111218 531922 111454
rect 531686 110898 531922 111134
rect 540686 111218 540922 111454
rect 540686 110898 540922 111134
rect 549686 111218 549922 111454
rect 549686 110898 549922 111134
rect 551488 111218 551724 111454
rect 551488 110898 551724 111134
rect 552860 111218 553096 111454
rect 552860 110898 553096 111134
rect 553706 111218 553942 111454
rect 553706 110898 553942 111134
rect 562706 111218 562942 111454
rect 562706 110898 562942 111134
rect 571706 111218 571942 111454
rect 571706 110898 571942 111134
rect 573476 111218 573712 111454
rect 573476 110898 573712 111134
rect 578670 111218 578906 111454
rect 578670 110898 578906 111134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 4582 93218 4818 93454
rect 4582 92898 4818 93134
rect 12232 93218 12468 93454
rect 12232 92898 12468 93134
rect 13038 93218 13274 93454
rect 13038 92898 13274 93134
rect 22038 93218 22274 93454
rect 22038 92898 22274 93134
rect 27588 93218 27824 93454
rect 27588 92898 27824 93134
rect 28240 93218 28476 93454
rect 28240 92898 28476 93134
rect 29046 93218 29282 93454
rect 29046 92898 29282 93134
rect 38046 93218 38282 93454
rect 38046 92898 38282 93134
rect 47046 93218 47282 93454
rect 47046 92898 47282 93134
rect 56046 93218 56282 93454
rect 56046 92898 56282 93134
rect 65046 93218 65282 93454
rect 65046 92898 65282 93134
rect 67608 93218 67844 93454
rect 67608 92898 67844 93134
rect 68260 93218 68496 93454
rect 68260 92898 68496 93134
rect 69066 93218 69302 93454
rect 69066 92898 69302 93134
rect 78066 93218 78302 93454
rect 78066 92898 78302 93134
rect 87066 93218 87302 93454
rect 87066 92898 87302 93134
rect 96066 93218 96302 93454
rect 96066 92898 96302 93134
rect 105066 93218 105302 93454
rect 105066 92898 105302 93134
rect 107628 93218 107864 93454
rect 107628 92898 107864 93134
rect 108280 93218 108516 93454
rect 108280 92898 108516 93134
rect 109086 93218 109322 93454
rect 109086 92898 109322 93134
rect 118086 93218 118322 93454
rect 118086 92898 118322 93134
rect 127086 93218 127322 93454
rect 127086 92898 127322 93134
rect 136086 93218 136322 93454
rect 136086 92898 136322 93134
rect 145086 93218 145322 93454
rect 145086 92898 145322 93134
rect 147648 93218 147884 93454
rect 147648 92898 147884 93134
rect 149300 93218 149536 93454
rect 149300 92898 149536 93134
rect 150106 93218 150342 93454
rect 150106 92898 150342 93134
rect 159106 93218 159342 93454
rect 159106 92898 159342 93134
rect 168106 93218 168342 93454
rect 168106 92898 168342 93134
rect 177106 93218 177342 93454
rect 177106 92898 177342 93134
rect 186106 93218 186342 93454
rect 186106 92898 186342 93134
rect 188668 93218 188904 93454
rect 188668 92898 188904 93134
rect 190320 93218 190556 93454
rect 190320 92898 190556 93134
rect 191126 93218 191362 93454
rect 191126 92898 191362 93134
rect 200126 93218 200362 93454
rect 200126 92898 200362 93134
rect 209126 93218 209362 93454
rect 209126 92898 209362 93134
rect 218126 93218 218362 93454
rect 218126 92898 218362 93134
rect 227126 93218 227362 93454
rect 227126 92898 227362 93134
rect 229688 93218 229924 93454
rect 229688 92898 229924 93134
rect 230340 93218 230576 93454
rect 230340 92898 230576 93134
rect 231146 93218 231382 93454
rect 231146 92898 231382 93134
rect 240146 93218 240382 93454
rect 240146 92898 240382 93134
rect 249146 93218 249382 93454
rect 249146 92898 249382 93134
rect 258146 93218 258382 93454
rect 258146 92898 258382 93134
rect 267146 93218 267382 93454
rect 267146 92898 267382 93134
rect 269708 93218 269944 93454
rect 269708 92898 269944 93134
rect 270360 93218 270596 93454
rect 270360 92898 270596 93134
rect 271166 93218 271402 93454
rect 271166 92898 271402 93134
rect 280166 93218 280402 93454
rect 280166 92898 280402 93134
rect 289166 93218 289402 93454
rect 289166 92898 289402 93134
rect 298166 93218 298402 93454
rect 298166 92898 298402 93134
rect 307166 93218 307402 93454
rect 307166 92898 307402 93134
rect 309728 93218 309964 93454
rect 309728 92898 309964 93134
rect 311380 93218 311616 93454
rect 311380 92898 311616 93134
rect 312186 93218 312422 93454
rect 312186 92898 312422 93134
rect 321186 93218 321422 93454
rect 321186 92898 321422 93134
rect 330186 93218 330422 93454
rect 330186 92898 330422 93134
rect 339186 93218 339422 93454
rect 339186 92898 339422 93134
rect 348186 93218 348422 93454
rect 348186 92898 348422 93134
rect 350748 93218 350984 93454
rect 350748 92898 350984 93134
rect 352400 93218 352636 93454
rect 352400 92898 352636 93134
rect 353206 93218 353442 93454
rect 353206 92898 353442 93134
rect 362206 93218 362442 93454
rect 362206 92898 362442 93134
rect 371206 93218 371442 93454
rect 371206 92898 371442 93134
rect 380206 93218 380442 93454
rect 380206 92898 380442 93134
rect 389206 93218 389442 93454
rect 389206 92898 389442 93134
rect 391768 93218 392004 93454
rect 391768 92898 392004 93134
rect 392420 93218 392656 93454
rect 392420 92898 392656 93134
rect 393226 93218 393462 93454
rect 393226 92898 393462 93134
rect 402226 93218 402462 93454
rect 402226 92898 402462 93134
rect 411226 93218 411462 93454
rect 411226 92898 411462 93134
rect 420226 93218 420462 93454
rect 420226 92898 420462 93134
rect 429226 93218 429462 93454
rect 429226 92898 429462 93134
rect 431788 93218 432024 93454
rect 431788 92898 432024 93134
rect 432440 93218 432676 93454
rect 432440 92898 432676 93134
rect 433246 93218 433482 93454
rect 433246 92898 433482 93134
rect 442246 93218 442482 93454
rect 442246 92898 442482 93134
rect 451246 93218 451482 93454
rect 451246 92898 451482 93134
rect 460246 93218 460482 93454
rect 460246 92898 460482 93134
rect 469246 93218 469482 93454
rect 469246 92898 469482 93134
rect 471808 93218 472044 93454
rect 471808 92898 472044 93134
rect 472460 93218 472696 93454
rect 472460 92898 472696 93134
rect 473266 93218 473502 93454
rect 473266 92898 473502 93134
rect 482266 93218 482502 93454
rect 482266 92898 482502 93134
rect 491266 93218 491502 93454
rect 491266 92898 491502 93134
rect 500266 93218 500502 93454
rect 500266 92898 500502 93134
rect 509266 93218 509502 93454
rect 509266 92898 509502 93134
rect 511828 93218 512064 93454
rect 511828 92898 512064 93134
rect 512480 93218 512716 93454
rect 512480 92898 512716 93134
rect 513286 93218 513522 93454
rect 513286 92898 513522 93134
rect 522286 93218 522522 93454
rect 522286 92898 522522 93134
rect 531286 93218 531522 93454
rect 531286 92898 531522 93134
rect 540286 93218 540522 93454
rect 540286 92898 540522 93134
rect 549286 93218 549522 93454
rect 549286 92898 549522 93134
rect 551848 93218 552084 93454
rect 551848 92898 552084 93134
rect 552500 93218 552736 93454
rect 552500 92898 552736 93134
rect 553306 93218 553542 93454
rect 553306 92898 553542 93134
rect 562306 93218 562542 93454
rect 562306 92898 562542 93134
rect 571306 93218 571542 93454
rect 571306 92898 571542 93134
rect 573836 93218 574072 93454
rect 573836 92898 574072 93134
rect 579470 93218 579706 93454
rect 579470 92898 579706 93134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect 5382 75218 5618 75454
rect 5382 74898 5618 75134
rect 12592 75218 12828 75454
rect 12592 74898 12828 75134
rect 13438 75218 13674 75454
rect 13438 74898 13674 75134
rect 22438 75218 22674 75454
rect 22438 74898 22674 75134
rect 27228 75218 27464 75454
rect 27228 74898 27464 75134
rect 28600 75218 28836 75454
rect 28600 74898 28836 75134
rect 29446 75218 29682 75454
rect 29446 74898 29682 75134
rect 38446 75218 38682 75454
rect 38446 74898 38682 75134
rect 47446 75218 47682 75454
rect 47446 74898 47682 75134
rect 56446 75218 56682 75454
rect 56446 74898 56682 75134
rect 65446 75218 65682 75454
rect 65446 74898 65682 75134
rect 67248 75218 67484 75454
rect 67248 74898 67484 75134
rect 68620 75218 68856 75454
rect 68620 74898 68856 75134
rect 69466 75218 69702 75454
rect 69466 74898 69702 75134
rect 78466 75218 78702 75454
rect 78466 74898 78702 75134
rect 87466 75218 87702 75454
rect 87466 74898 87702 75134
rect 96466 75218 96702 75454
rect 96466 74898 96702 75134
rect 105466 75218 105702 75454
rect 105466 74898 105702 75134
rect 107268 75218 107504 75454
rect 107268 74898 107504 75134
rect 108640 75218 108876 75454
rect 108640 74898 108876 75134
rect 109486 75218 109722 75454
rect 109486 74898 109722 75134
rect 118486 75218 118722 75454
rect 118486 74898 118722 75134
rect 127486 75218 127722 75454
rect 127486 74898 127722 75134
rect 136486 75218 136722 75454
rect 136486 74898 136722 75134
rect 145486 75218 145722 75454
rect 145486 74898 145722 75134
rect 147288 75218 147524 75454
rect 147288 74898 147524 75134
rect 149660 75218 149896 75454
rect 149660 74898 149896 75134
rect 150506 75218 150742 75454
rect 150506 74898 150742 75134
rect 159506 75218 159742 75454
rect 159506 74898 159742 75134
rect 168506 75218 168742 75454
rect 168506 74898 168742 75134
rect 177506 75218 177742 75454
rect 177506 74898 177742 75134
rect 186506 75218 186742 75454
rect 186506 74898 186742 75134
rect 188308 75218 188544 75454
rect 188308 74898 188544 75134
rect 190680 75218 190916 75454
rect 190680 74898 190916 75134
rect 191526 75218 191762 75454
rect 191526 74898 191762 75134
rect 200526 75218 200762 75454
rect 200526 74898 200762 75134
rect 209526 75218 209762 75454
rect 209526 74898 209762 75134
rect 218526 75218 218762 75454
rect 218526 74898 218762 75134
rect 227526 75218 227762 75454
rect 227526 74898 227762 75134
rect 229328 75218 229564 75454
rect 229328 74898 229564 75134
rect 230700 75218 230936 75454
rect 230700 74898 230936 75134
rect 231546 75218 231782 75454
rect 231546 74898 231782 75134
rect 240546 75218 240782 75454
rect 240546 74898 240782 75134
rect 249546 75218 249782 75454
rect 249546 74898 249782 75134
rect 258546 75218 258782 75454
rect 258546 74898 258782 75134
rect 267546 75218 267782 75454
rect 267546 74898 267782 75134
rect 269348 75218 269584 75454
rect 269348 74898 269584 75134
rect 270720 75218 270956 75454
rect 270720 74898 270956 75134
rect 271566 75218 271802 75454
rect 271566 74898 271802 75134
rect 280566 75218 280802 75454
rect 280566 74898 280802 75134
rect 289566 75218 289802 75454
rect 289566 74898 289802 75134
rect 298566 75218 298802 75454
rect 298566 74898 298802 75134
rect 307566 75218 307802 75454
rect 307566 74898 307802 75134
rect 309368 75218 309604 75454
rect 309368 74898 309604 75134
rect 311740 75218 311976 75454
rect 311740 74898 311976 75134
rect 312586 75218 312822 75454
rect 312586 74898 312822 75134
rect 321586 75218 321822 75454
rect 321586 74898 321822 75134
rect 330586 75218 330822 75454
rect 330586 74898 330822 75134
rect 339586 75218 339822 75454
rect 339586 74898 339822 75134
rect 348586 75218 348822 75454
rect 348586 74898 348822 75134
rect 350388 75218 350624 75454
rect 350388 74898 350624 75134
rect 352760 75218 352996 75454
rect 352760 74898 352996 75134
rect 353606 75218 353842 75454
rect 353606 74898 353842 75134
rect 362606 75218 362842 75454
rect 362606 74898 362842 75134
rect 371606 75218 371842 75454
rect 371606 74898 371842 75134
rect 380606 75218 380842 75454
rect 380606 74898 380842 75134
rect 389606 75218 389842 75454
rect 389606 74898 389842 75134
rect 391408 75218 391644 75454
rect 391408 74898 391644 75134
rect 392780 75218 393016 75454
rect 392780 74898 393016 75134
rect 393626 75218 393862 75454
rect 393626 74898 393862 75134
rect 402626 75218 402862 75454
rect 402626 74898 402862 75134
rect 411626 75218 411862 75454
rect 411626 74898 411862 75134
rect 420626 75218 420862 75454
rect 420626 74898 420862 75134
rect 429626 75218 429862 75454
rect 429626 74898 429862 75134
rect 431428 75218 431664 75454
rect 431428 74898 431664 75134
rect 432800 75218 433036 75454
rect 432800 74898 433036 75134
rect 433646 75218 433882 75454
rect 433646 74898 433882 75134
rect 442646 75218 442882 75454
rect 442646 74898 442882 75134
rect 451646 75218 451882 75454
rect 451646 74898 451882 75134
rect 460646 75218 460882 75454
rect 460646 74898 460882 75134
rect 469646 75218 469882 75454
rect 469646 74898 469882 75134
rect 471448 75218 471684 75454
rect 471448 74898 471684 75134
rect 472820 75218 473056 75454
rect 472820 74898 473056 75134
rect 473666 75218 473902 75454
rect 473666 74898 473902 75134
rect 482666 75218 482902 75454
rect 482666 74898 482902 75134
rect 491666 75218 491902 75454
rect 491666 74898 491902 75134
rect 500666 75218 500902 75454
rect 500666 74898 500902 75134
rect 509666 75218 509902 75454
rect 509666 74898 509902 75134
rect 511468 75218 511704 75454
rect 511468 74898 511704 75134
rect 512840 75218 513076 75454
rect 512840 74898 513076 75134
rect 513686 75218 513922 75454
rect 513686 74898 513922 75134
rect 522686 75218 522922 75454
rect 522686 74898 522922 75134
rect 531686 75218 531922 75454
rect 531686 74898 531922 75134
rect 540686 75218 540922 75454
rect 540686 74898 540922 75134
rect 549686 75218 549922 75454
rect 549686 74898 549922 75134
rect 551488 75218 551724 75454
rect 551488 74898 551724 75134
rect 552860 75218 553096 75454
rect 552860 74898 553096 75134
rect 553706 75218 553942 75454
rect 553706 74898 553942 75134
rect 562706 75218 562942 75454
rect 562706 74898 562942 75134
rect 571706 75218 571942 75454
rect 571706 74898 571942 75134
rect 573476 75218 573712 75454
rect 573476 74898 573712 75134
rect 578670 75218 578906 75454
rect 578670 74898 578906 75134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 4582 57218 4818 57454
rect 4582 56898 4818 57134
rect 28240 57218 28476 57454
rect 28240 56898 28476 57134
rect 29046 57218 29282 57454
rect 29046 56898 29282 57134
rect 38046 57218 38282 57454
rect 38046 56898 38282 57134
rect 47046 57218 47282 57454
rect 47046 56898 47282 57134
rect 56046 57218 56282 57454
rect 56046 56898 56282 57134
rect 65046 57218 65282 57454
rect 65046 56898 65282 57134
rect 67608 57218 67844 57454
rect 67608 56898 67844 57134
rect 68260 57218 68496 57454
rect 68260 56898 68496 57134
rect 69066 57218 69302 57454
rect 69066 56898 69302 57134
rect 78066 57218 78302 57454
rect 78066 56898 78302 57134
rect 87066 57218 87302 57454
rect 87066 56898 87302 57134
rect 96066 57218 96302 57454
rect 96066 56898 96302 57134
rect 105066 57218 105302 57454
rect 105066 56898 105302 57134
rect 107628 57218 107864 57454
rect 107628 56898 107864 57134
rect 108280 57218 108516 57454
rect 108280 56898 108516 57134
rect 109086 57218 109322 57454
rect 109086 56898 109322 57134
rect 118086 57218 118322 57454
rect 118086 56898 118322 57134
rect 127086 57218 127322 57454
rect 127086 56898 127322 57134
rect 136086 57218 136322 57454
rect 136086 56898 136322 57134
rect 145086 57218 145322 57454
rect 145086 56898 145322 57134
rect 147648 57218 147884 57454
rect 147648 56898 147884 57134
rect 149300 57218 149536 57454
rect 149300 56898 149536 57134
rect 150106 57218 150342 57454
rect 150106 56898 150342 57134
rect 159106 57218 159342 57454
rect 159106 56898 159342 57134
rect 168106 57218 168342 57454
rect 168106 56898 168342 57134
rect 177106 57218 177342 57454
rect 177106 56898 177342 57134
rect 186106 57218 186342 57454
rect 186106 56898 186342 57134
rect 188668 57218 188904 57454
rect 188668 56898 188904 57134
rect 190320 57218 190556 57454
rect 190320 56898 190556 57134
rect 191126 57218 191362 57454
rect 191126 56898 191362 57134
rect 200126 57218 200362 57454
rect 200126 56898 200362 57134
rect 209126 57218 209362 57454
rect 209126 56898 209362 57134
rect 218126 57218 218362 57454
rect 218126 56898 218362 57134
rect 227126 57218 227362 57454
rect 227126 56898 227362 57134
rect 229688 57218 229924 57454
rect 229688 56898 229924 57134
rect 230340 57218 230576 57454
rect 230340 56898 230576 57134
rect 231146 57218 231382 57454
rect 231146 56898 231382 57134
rect 240146 57218 240382 57454
rect 240146 56898 240382 57134
rect 249146 57218 249382 57454
rect 249146 56898 249382 57134
rect 258146 57218 258382 57454
rect 258146 56898 258382 57134
rect 267146 57218 267382 57454
rect 267146 56898 267382 57134
rect 269708 57218 269944 57454
rect 269708 56898 269944 57134
rect 270360 57218 270596 57454
rect 270360 56898 270596 57134
rect 271166 57218 271402 57454
rect 271166 56898 271402 57134
rect 280166 57218 280402 57454
rect 280166 56898 280402 57134
rect 289166 57218 289402 57454
rect 289166 56898 289402 57134
rect 298166 57218 298402 57454
rect 298166 56898 298402 57134
rect 307166 57218 307402 57454
rect 307166 56898 307402 57134
rect 309728 57218 309964 57454
rect 309728 56898 309964 57134
rect 311380 57218 311616 57454
rect 311380 56898 311616 57134
rect 312186 57218 312422 57454
rect 312186 56898 312422 57134
rect 321186 57218 321422 57454
rect 321186 56898 321422 57134
rect 330186 57218 330422 57454
rect 330186 56898 330422 57134
rect 339186 57218 339422 57454
rect 339186 56898 339422 57134
rect 348186 57218 348422 57454
rect 348186 56898 348422 57134
rect 350748 57218 350984 57454
rect 350748 56898 350984 57134
rect 352400 57218 352636 57454
rect 352400 56898 352636 57134
rect 353206 57218 353442 57454
rect 353206 56898 353442 57134
rect 362206 57218 362442 57454
rect 362206 56898 362442 57134
rect 371206 57218 371442 57454
rect 371206 56898 371442 57134
rect 380206 57218 380442 57454
rect 380206 56898 380442 57134
rect 389206 57218 389442 57454
rect 389206 56898 389442 57134
rect 391768 57218 392004 57454
rect 391768 56898 392004 57134
rect 392420 57218 392656 57454
rect 392420 56898 392656 57134
rect 393226 57218 393462 57454
rect 393226 56898 393462 57134
rect 402226 57218 402462 57454
rect 402226 56898 402462 57134
rect 411226 57218 411462 57454
rect 411226 56898 411462 57134
rect 420226 57218 420462 57454
rect 420226 56898 420462 57134
rect 429226 57218 429462 57454
rect 429226 56898 429462 57134
rect 431788 57218 432024 57454
rect 431788 56898 432024 57134
rect 432440 57218 432676 57454
rect 432440 56898 432676 57134
rect 433246 57218 433482 57454
rect 433246 56898 433482 57134
rect 442246 57218 442482 57454
rect 442246 56898 442482 57134
rect 451246 57218 451482 57454
rect 451246 56898 451482 57134
rect 460246 57218 460482 57454
rect 460246 56898 460482 57134
rect 469246 57218 469482 57454
rect 469246 56898 469482 57134
rect 471808 57218 472044 57454
rect 471808 56898 472044 57134
rect 472460 57218 472696 57454
rect 472460 56898 472696 57134
rect 473266 57218 473502 57454
rect 473266 56898 473502 57134
rect 482266 57218 482502 57454
rect 482266 56898 482502 57134
rect 491266 57218 491502 57454
rect 491266 56898 491502 57134
rect 500266 57218 500502 57454
rect 500266 56898 500502 57134
rect 509266 57218 509502 57454
rect 509266 56898 509502 57134
rect 511828 57218 512064 57454
rect 511828 56898 512064 57134
rect 512480 57218 512716 57454
rect 512480 56898 512716 57134
rect 513286 57218 513522 57454
rect 513286 56898 513522 57134
rect 522286 57218 522522 57454
rect 522286 56898 522522 57134
rect 531286 57218 531522 57454
rect 531286 56898 531522 57134
rect 540286 57218 540522 57454
rect 540286 56898 540522 57134
rect 549286 57218 549522 57454
rect 549286 56898 549522 57134
rect 551848 57218 552084 57454
rect 551848 56898 552084 57134
rect 552500 57218 552736 57454
rect 552500 56898 552736 57134
rect 553306 57218 553542 57454
rect 553306 56898 553542 57134
rect 562306 57218 562542 57454
rect 562306 56898 562542 57134
rect 571306 57218 571542 57454
rect 571306 56898 571542 57134
rect 573836 57218 574072 57454
rect 573836 56898 574072 57134
rect 579470 57218 579706 57454
rect 579470 56898 579706 57134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect 5382 39218 5618 39454
rect 5382 38898 5618 39134
rect 578670 39218 578906 39454
rect 578670 38898 578906 39134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 4582 669454
rect 4818 669218 127058 669454
rect 127294 669218 140296 669454
rect 140532 669218 147648 669454
rect 147884 669218 190320 669454
rect 190556 669218 229688 669454
rect 229924 669218 432440 669454
rect 432676 669218 439792 669454
rect 440028 669218 457010 669454
rect 457246 669218 579470 669454
rect 579706 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 4582 669134
rect 4818 668898 127058 669134
rect 127294 668898 140296 669134
rect 140532 668898 147648 669134
rect 147884 668898 190320 669134
rect 190556 668898 229688 669134
rect 229924 668898 432440 669134
rect 432676 668898 439792 669134
rect 440028 668898 457010 669134
rect 457246 668898 579470 669134
rect 579706 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 5382 651454
rect 5618 651218 127458 651454
rect 127694 651218 140656 651454
rect 140892 651218 147288 651454
rect 147524 651218 149660 651454
rect 149896 651218 188308 651454
rect 188544 651218 190680 651454
rect 190916 651218 229328 651454
rect 229564 651218 230700 651454
rect 230936 651218 269348 651454
rect 269584 651218 270720 651454
rect 270956 651218 309368 651454
rect 309604 651218 310564 651454
rect 310800 651218 311740 651454
rect 311976 651218 350388 651454
rect 350624 651218 352760 651454
rect 352996 651218 391408 651454
rect 391644 651218 392780 651454
rect 393016 651218 431428 651454
rect 431664 651218 432800 651454
rect 433036 651218 439432 651454
rect 439668 651218 456610 651454
rect 456846 651218 578670 651454
rect 578906 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 5382 651134
rect 5618 650898 127458 651134
rect 127694 650898 140656 651134
rect 140892 650898 147288 651134
rect 147524 650898 149660 651134
rect 149896 650898 188308 651134
rect 188544 650898 190680 651134
rect 190916 650898 229328 651134
rect 229564 650898 230700 651134
rect 230936 650898 269348 651134
rect 269584 650898 270720 651134
rect 270956 650898 309368 651134
rect 309604 650898 310564 651134
rect 310800 650898 311740 651134
rect 311976 650898 350388 651134
rect 350624 650898 352760 651134
rect 352996 650898 391408 651134
rect 391644 650898 392780 651134
rect 393016 650898 431428 651134
rect 431664 650898 432800 651134
rect 433036 650898 439432 651134
rect 439668 650898 456610 651134
rect 456846 650898 578670 651134
rect 578906 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 4582 633454
rect 4818 633218 12352 633454
rect 12588 633218 107416 633454
rect 107652 633218 127058 633454
rect 127294 633218 140296 633454
rect 140532 633218 141102 633454
rect 141338 633218 147648 633454
rect 147884 633218 149300 633454
rect 149536 633218 150106 633454
rect 150342 633218 159106 633454
rect 159342 633218 168106 633454
rect 168342 633218 177106 633454
rect 177342 633218 186106 633454
rect 186342 633218 188668 633454
rect 188904 633218 190320 633454
rect 190556 633218 191126 633454
rect 191362 633218 200126 633454
rect 200362 633218 209126 633454
rect 209362 633218 218126 633454
rect 218362 633218 227126 633454
rect 227362 633218 229688 633454
rect 229924 633218 230340 633454
rect 230576 633218 231146 633454
rect 231382 633218 240146 633454
rect 240382 633218 249146 633454
rect 249382 633218 258146 633454
rect 258382 633218 267146 633454
rect 267382 633218 269708 633454
rect 269944 633218 270360 633454
rect 270596 633218 271166 633454
rect 271402 633218 280166 633454
rect 280402 633218 289166 633454
rect 289402 633218 298166 633454
rect 298402 633218 307166 633454
rect 307402 633218 309728 633454
rect 309964 633218 311380 633454
rect 311616 633218 312186 633454
rect 312422 633218 321186 633454
rect 321422 633218 330186 633454
rect 330422 633218 339186 633454
rect 339422 633218 348186 633454
rect 348422 633218 350748 633454
rect 350984 633218 352400 633454
rect 352636 633218 353206 633454
rect 353442 633218 362206 633454
rect 362442 633218 371206 633454
rect 371442 633218 380206 633454
rect 380442 633218 389206 633454
rect 389442 633218 391768 633454
rect 392004 633218 392420 633454
rect 392656 633218 393226 633454
rect 393462 633218 402226 633454
rect 402462 633218 411226 633454
rect 411462 633218 420226 633454
rect 420462 633218 429226 633454
rect 429462 633218 431788 633454
rect 432024 633218 432440 633454
rect 432676 633218 433246 633454
rect 433482 633218 439792 633454
rect 440028 633218 457010 633454
rect 457246 633218 476652 633454
rect 476888 633218 571716 633454
rect 571952 633218 579470 633454
rect 579706 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 4582 633134
rect 4818 632898 12352 633134
rect 12588 632898 107416 633134
rect 107652 632898 127058 633134
rect 127294 632898 140296 633134
rect 140532 632898 141102 633134
rect 141338 632898 147648 633134
rect 147884 632898 149300 633134
rect 149536 632898 150106 633134
rect 150342 632898 159106 633134
rect 159342 632898 168106 633134
rect 168342 632898 177106 633134
rect 177342 632898 186106 633134
rect 186342 632898 188668 633134
rect 188904 632898 190320 633134
rect 190556 632898 191126 633134
rect 191362 632898 200126 633134
rect 200362 632898 209126 633134
rect 209362 632898 218126 633134
rect 218362 632898 227126 633134
rect 227362 632898 229688 633134
rect 229924 632898 230340 633134
rect 230576 632898 231146 633134
rect 231382 632898 240146 633134
rect 240382 632898 249146 633134
rect 249382 632898 258146 633134
rect 258382 632898 267146 633134
rect 267382 632898 269708 633134
rect 269944 632898 270360 633134
rect 270596 632898 271166 633134
rect 271402 632898 280166 633134
rect 280402 632898 289166 633134
rect 289402 632898 298166 633134
rect 298402 632898 307166 633134
rect 307402 632898 309728 633134
rect 309964 632898 311380 633134
rect 311616 632898 312186 633134
rect 312422 632898 321186 633134
rect 321422 632898 330186 633134
rect 330422 632898 339186 633134
rect 339422 632898 348186 633134
rect 348422 632898 350748 633134
rect 350984 632898 352400 633134
rect 352636 632898 353206 633134
rect 353442 632898 362206 633134
rect 362442 632898 371206 633134
rect 371442 632898 380206 633134
rect 380442 632898 389206 633134
rect 389442 632898 391768 633134
rect 392004 632898 392420 633134
rect 392656 632898 393226 633134
rect 393462 632898 402226 633134
rect 402462 632898 411226 633134
rect 411462 632898 420226 633134
rect 420462 632898 429226 633134
rect 429462 632898 431788 633134
rect 432024 632898 432440 633134
rect 432676 632898 433246 633134
rect 433482 632898 439792 633134
rect 440028 632898 457010 633134
rect 457246 632898 476652 633134
rect 476888 632898 571716 633134
rect 571952 632898 579470 633134
rect 579706 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 5382 615454
rect 5618 615218 13032 615454
rect 13268 615218 106736 615454
rect 106972 615218 127458 615454
rect 127694 615218 140656 615454
rect 140892 615218 141502 615454
rect 141738 615218 147288 615454
rect 147524 615218 149660 615454
rect 149896 615218 150506 615454
rect 150742 615218 159506 615454
rect 159742 615218 168506 615454
rect 168742 615218 177506 615454
rect 177742 615218 186506 615454
rect 186742 615218 188308 615454
rect 188544 615218 190680 615454
rect 190916 615218 191526 615454
rect 191762 615218 200526 615454
rect 200762 615218 209526 615454
rect 209762 615218 218526 615454
rect 218762 615218 227526 615454
rect 227762 615218 229328 615454
rect 229564 615218 230700 615454
rect 230936 615218 231546 615454
rect 231782 615218 240546 615454
rect 240782 615218 249546 615454
rect 249782 615218 258546 615454
rect 258782 615218 267546 615454
rect 267782 615218 269348 615454
rect 269584 615218 270720 615454
rect 270956 615218 271566 615454
rect 271802 615218 280566 615454
rect 280802 615218 289566 615454
rect 289802 615218 298566 615454
rect 298802 615218 307566 615454
rect 307802 615218 309368 615454
rect 309604 615218 311740 615454
rect 311976 615218 312586 615454
rect 312822 615218 321586 615454
rect 321822 615218 330586 615454
rect 330822 615218 339586 615454
rect 339822 615218 348586 615454
rect 348822 615218 350388 615454
rect 350624 615218 352760 615454
rect 352996 615218 353606 615454
rect 353842 615218 362606 615454
rect 362842 615218 371606 615454
rect 371842 615218 380606 615454
rect 380842 615218 389606 615454
rect 389842 615218 391408 615454
rect 391644 615218 392780 615454
rect 393016 615218 393626 615454
rect 393862 615218 402626 615454
rect 402862 615218 411626 615454
rect 411862 615218 420626 615454
rect 420862 615218 429626 615454
rect 429862 615218 431428 615454
rect 431664 615218 432800 615454
rect 433036 615218 433646 615454
rect 433882 615218 439432 615454
rect 439668 615218 456610 615454
rect 456846 615218 477332 615454
rect 477568 615218 571036 615454
rect 571272 615218 578670 615454
rect 578906 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 5382 615134
rect 5618 614898 13032 615134
rect 13268 614898 106736 615134
rect 106972 614898 127458 615134
rect 127694 614898 140656 615134
rect 140892 614898 141502 615134
rect 141738 614898 147288 615134
rect 147524 614898 149660 615134
rect 149896 614898 150506 615134
rect 150742 614898 159506 615134
rect 159742 614898 168506 615134
rect 168742 614898 177506 615134
rect 177742 614898 186506 615134
rect 186742 614898 188308 615134
rect 188544 614898 190680 615134
rect 190916 614898 191526 615134
rect 191762 614898 200526 615134
rect 200762 614898 209526 615134
rect 209762 614898 218526 615134
rect 218762 614898 227526 615134
rect 227762 614898 229328 615134
rect 229564 614898 230700 615134
rect 230936 614898 231546 615134
rect 231782 614898 240546 615134
rect 240782 614898 249546 615134
rect 249782 614898 258546 615134
rect 258782 614898 267546 615134
rect 267782 614898 269348 615134
rect 269584 614898 270720 615134
rect 270956 614898 271566 615134
rect 271802 614898 280566 615134
rect 280802 614898 289566 615134
rect 289802 614898 298566 615134
rect 298802 614898 307566 615134
rect 307802 614898 309368 615134
rect 309604 614898 311740 615134
rect 311976 614898 312586 615134
rect 312822 614898 321586 615134
rect 321822 614898 330586 615134
rect 330822 614898 339586 615134
rect 339822 614898 348586 615134
rect 348822 614898 350388 615134
rect 350624 614898 352760 615134
rect 352996 614898 353606 615134
rect 353842 614898 362606 615134
rect 362842 614898 371606 615134
rect 371842 614898 380606 615134
rect 380842 614898 389606 615134
rect 389842 614898 391408 615134
rect 391644 614898 392780 615134
rect 393016 614898 393626 615134
rect 393862 614898 402626 615134
rect 402862 614898 411626 615134
rect 411862 614898 420626 615134
rect 420862 614898 429626 615134
rect 429862 614898 431428 615134
rect 431664 614898 432800 615134
rect 433036 614898 433646 615134
rect 433882 614898 439432 615134
rect 439668 614898 456610 615134
rect 456846 614898 477332 615134
rect 477568 614898 571036 615134
rect 571272 614898 578670 615134
rect 578906 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 4582 597454
rect 4818 597218 12352 597454
rect 12588 597218 107416 597454
rect 107652 597218 127058 597454
rect 127294 597218 140296 597454
rect 140532 597218 141102 597454
rect 141338 597218 147648 597454
rect 147884 597218 149300 597454
rect 149536 597218 150106 597454
rect 150342 597218 159106 597454
rect 159342 597218 168106 597454
rect 168342 597218 177106 597454
rect 177342 597218 186106 597454
rect 186342 597218 188668 597454
rect 188904 597218 189768 597454
rect 190004 597218 190320 597454
rect 190556 597218 191126 597454
rect 191362 597218 200126 597454
rect 200362 597218 209126 597454
rect 209362 597218 218126 597454
rect 218362 597218 227126 597454
rect 227362 597218 229688 597454
rect 229924 597218 230340 597454
rect 230576 597218 231146 597454
rect 231382 597218 240146 597454
rect 240382 597218 249146 597454
rect 249382 597218 258146 597454
rect 258382 597218 267146 597454
rect 267382 597218 269708 597454
rect 269944 597218 270360 597454
rect 270596 597218 271166 597454
rect 271402 597218 280166 597454
rect 280402 597218 289166 597454
rect 289402 597218 298166 597454
rect 298402 597218 307166 597454
rect 307402 597218 309728 597454
rect 309964 597218 311380 597454
rect 311616 597218 312186 597454
rect 312422 597218 321186 597454
rect 321422 597218 330186 597454
rect 330422 597218 339186 597454
rect 339422 597218 348186 597454
rect 348422 597218 350748 597454
rect 350984 597218 352400 597454
rect 352636 597218 353206 597454
rect 353442 597218 362206 597454
rect 362442 597218 371206 597454
rect 371442 597218 380206 597454
rect 380442 597218 389206 597454
rect 389442 597218 391768 597454
rect 392004 597218 392420 597454
rect 392656 597218 393226 597454
rect 393462 597218 402226 597454
rect 402462 597218 411226 597454
rect 411462 597218 420226 597454
rect 420462 597218 429226 597454
rect 429462 597218 431788 597454
rect 432024 597218 432440 597454
rect 432676 597218 433246 597454
rect 433482 597218 439792 597454
rect 440028 597218 457010 597454
rect 457246 597218 476652 597454
rect 476888 597218 571716 597454
rect 571952 597218 579470 597454
rect 579706 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 4582 597134
rect 4818 596898 12352 597134
rect 12588 596898 107416 597134
rect 107652 596898 127058 597134
rect 127294 596898 140296 597134
rect 140532 596898 141102 597134
rect 141338 596898 147648 597134
rect 147884 596898 149300 597134
rect 149536 596898 150106 597134
rect 150342 596898 159106 597134
rect 159342 596898 168106 597134
rect 168342 596898 177106 597134
rect 177342 596898 186106 597134
rect 186342 596898 188668 597134
rect 188904 596898 189768 597134
rect 190004 596898 190320 597134
rect 190556 596898 191126 597134
rect 191362 596898 200126 597134
rect 200362 596898 209126 597134
rect 209362 596898 218126 597134
rect 218362 596898 227126 597134
rect 227362 596898 229688 597134
rect 229924 596898 230340 597134
rect 230576 596898 231146 597134
rect 231382 596898 240146 597134
rect 240382 596898 249146 597134
rect 249382 596898 258146 597134
rect 258382 596898 267146 597134
rect 267382 596898 269708 597134
rect 269944 596898 270360 597134
rect 270596 596898 271166 597134
rect 271402 596898 280166 597134
rect 280402 596898 289166 597134
rect 289402 596898 298166 597134
rect 298402 596898 307166 597134
rect 307402 596898 309728 597134
rect 309964 596898 311380 597134
rect 311616 596898 312186 597134
rect 312422 596898 321186 597134
rect 321422 596898 330186 597134
rect 330422 596898 339186 597134
rect 339422 596898 348186 597134
rect 348422 596898 350748 597134
rect 350984 596898 352400 597134
rect 352636 596898 353206 597134
rect 353442 596898 362206 597134
rect 362442 596898 371206 597134
rect 371442 596898 380206 597134
rect 380442 596898 389206 597134
rect 389442 596898 391768 597134
rect 392004 596898 392420 597134
rect 392656 596898 393226 597134
rect 393462 596898 402226 597134
rect 402462 596898 411226 597134
rect 411462 596898 420226 597134
rect 420462 596898 429226 597134
rect 429462 596898 431788 597134
rect 432024 596898 432440 597134
rect 432676 596898 433246 597134
rect 433482 596898 439792 597134
rect 440028 596898 457010 597134
rect 457246 596898 476652 597134
rect 476888 596898 571716 597134
rect 571952 596898 579470 597134
rect 579706 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 5382 579454
rect 5618 579218 13032 579454
rect 13268 579218 106736 579454
rect 106972 579218 127458 579454
rect 127694 579218 140656 579454
rect 140892 579218 141502 579454
rect 141738 579218 147288 579454
rect 147524 579218 149660 579454
rect 149896 579218 150506 579454
rect 150742 579218 159506 579454
rect 159742 579218 168506 579454
rect 168742 579218 177506 579454
rect 177742 579218 186506 579454
rect 186742 579218 188308 579454
rect 188544 579218 190680 579454
rect 190916 579218 191526 579454
rect 191762 579218 200526 579454
rect 200762 579218 209526 579454
rect 209762 579218 218526 579454
rect 218762 579218 227526 579454
rect 227762 579218 229328 579454
rect 229564 579218 230700 579454
rect 230936 579218 231546 579454
rect 231782 579218 240546 579454
rect 240782 579218 249546 579454
rect 249782 579218 258546 579454
rect 258782 579218 267546 579454
rect 267782 579218 269348 579454
rect 269584 579218 270720 579454
rect 270956 579218 271566 579454
rect 271802 579218 280566 579454
rect 280802 579218 289566 579454
rect 289802 579218 298566 579454
rect 298802 579218 307566 579454
rect 307802 579218 309368 579454
rect 309604 579218 311740 579454
rect 311976 579218 312586 579454
rect 312822 579218 321586 579454
rect 321822 579218 330586 579454
rect 330822 579218 339586 579454
rect 339822 579218 348586 579454
rect 348822 579218 350388 579454
rect 350624 579218 352760 579454
rect 352996 579218 353606 579454
rect 353842 579218 362606 579454
rect 362842 579218 371606 579454
rect 371842 579218 380606 579454
rect 380842 579218 389606 579454
rect 389842 579218 391408 579454
rect 391644 579218 392780 579454
rect 393016 579218 393626 579454
rect 393862 579218 402626 579454
rect 402862 579218 411626 579454
rect 411862 579218 420626 579454
rect 420862 579218 429626 579454
rect 429862 579218 431428 579454
rect 431664 579218 432800 579454
rect 433036 579218 433646 579454
rect 433882 579218 439432 579454
rect 439668 579218 456610 579454
rect 456846 579218 477332 579454
rect 477568 579218 571036 579454
rect 571272 579218 578670 579454
rect 578906 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 5382 579134
rect 5618 578898 13032 579134
rect 13268 578898 106736 579134
rect 106972 578898 127458 579134
rect 127694 578898 140656 579134
rect 140892 578898 141502 579134
rect 141738 578898 147288 579134
rect 147524 578898 149660 579134
rect 149896 578898 150506 579134
rect 150742 578898 159506 579134
rect 159742 578898 168506 579134
rect 168742 578898 177506 579134
rect 177742 578898 186506 579134
rect 186742 578898 188308 579134
rect 188544 578898 190680 579134
rect 190916 578898 191526 579134
rect 191762 578898 200526 579134
rect 200762 578898 209526 579134
rect 209762 578898 218526 579134
rect 218762 578898 227526 579134
rect 227762 578898 229328 579134
rect 229564 578898 230700 579134
rect 230936 578898 231546 579134
rect 231782 578898 240546 579134
rect 240782 578898 249546 579134
rect 249782 578898 258546 579134
rect 258782 578898 267546 579134
rect 267782 578898 269348 579134
rect 269584 578898 270720 579134
rect 270956 578898 271566 579134
rect 271802 578898 280566 579134
rect 280802 578898 289566 579134
rect 289802 578898 298566 579134
rect 298802 578898 307566 579134
rect 307802 578898 309368 579134
rect 309604 578898 311740 579134
rect 311976 578898 312586 579134
rect 312822 578898 321586 579134
rect 321822 578898 330586 579134
rect 330822 578898 339586 579134
rect 339822 578898 348586 579134
rect 348822 578898 350388 579134
rect 350624 578898 352760 579134
rect 352996 578898 353606 579134
rect 353842 578898 362606 579134
rect 362842 578898 371606 579134
rect 371842 578898 380606 579134
rect 380842 578898 389606 579134
rect 389842 578898 391408 579134
rect 391644 578898 392780 579134
rect 393016 578898 393626 579134
rect 393862 578898 402626 579134
rect 402862 578898 411626 579134
rect 411862 578898 420626 579134
rect 420862 578898 429626 579134
rect 429862 578898 431428 579134
rect 431664 578898 432800 579134
rect 433036 578898 433646 579134
rect 433882 578898 439432 579134
rect 439668 578898 456610 579134
rect 456846 578898 477332 579134
rect 477568 578898 571036 579134
rect 571272 578898 578670 579134
rect 578906 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 4582 561454
rect 4818 561218 12352 561454
rect 12588 561218 107416 561454
rect 107652 561218 127058 561454
rect 127294 561218 140296 561454
rect 140532 561218 141102 561454
rect 141338 561218 147648 561454
rect 147884 561218 149300 561454
rect 149536 561218 150106 561454
rect 150342 561218 159106 561454
rect 159342 561218 168106 561454
rect 168342 561218 177106 561454
rect 177342 561218 186106 561454
rect 186342 561218 188668 561454
rect 188904 561218 190320 561454
rect 190556 561218 191126 561454
rect 191362 561218 200126 561454
rect 200362 561218 209126 561454
rect 209362 561218 218126 561454
rect 218362 561218 227126 561454
rect 227362 561218 229688 561454
rect 229924 561218 230340 561454
rect 230576 561218 231146 561454
rect 231382 561218 240146 561454
rect 240382 561218 249146 561454
rect 249382 561218 258146 561454
rect 258382 561218 267146 561454
rect 267382 561218 269708 561454
rect 269944 561218 270360 561454
rect 270596 561218 271166 561454
rect 271402 561218 280166 561454
rect 280402 561218 289166 561454
rect 289402 561218 298166 561454
rect 298402 561218 307166 561454
rect 307402 561218 309728 561454
rect 309964 561218 311380 561454
rect 311616 561218 312186 561454
rect 312422 561218 321186 561454
rect 321422 561218 330186 561454
rect 330422 561218 339186 561454
rect 339422 561218 348186 561454
rect 348422 561218 350748 561454
rect 350984 561218 352400 561454
rect 352636 561218 353206 561454
rect 353442 561218 362206 561454
rect 362442 561218 371206 561454
rect 371442 561218 380206 561454
rect 380442 561218 389206 561454
rect 389442 561218 391768 561454
rect 392004 561218 392420 561454
rect 392656 561218 393226 561454
rect 393462 561218 402226 561454
rect 402462 561218 411226 561454
rect 411462 561218 420226 561454
rect 420462 561218 429226 561454
rect 429462 561218 431788 561454
rect 432024 561218 432440 561454
rect 432676 561218 433246 561454
rect 433482 561218 439792 561454
rect 440028 561218 457010 561454
rect 457246 561218 476652 561454
rect 476888 561218 571716 561454
rect 571952 561218 579470 561454
rect 579706 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 4582 561134
rect 4818 560898 12352 561134
rect 12588 560898 107416 561134
rect 107652 560898 127058 561134
rect 127294 560898 140296 561134
rect 140532 560898 141102 561134
rect 141338 560898 147648 561134
rect 147884 560898 149300 561134
rect 149536 560898 150106 561134
rect 150342 560898 159106 561134
rect 159342 560898 168106 561134
rect 168342 560898 177106 561134
rect 177342 560898 186106 561134
rect 186342 560898 188668 561134
rect 188904 560898 190320 561134
rect 190556 560898 191126 561134
rect 191362 560898 200126 561134
rect 200362 560898 209126 561134
rect 209362 560898 218126 561134
rect 218362 560898 227126 561134
rect 227362 560898 229688 561134
rect 229924 560898 230340 561134
rect 230576 560898 231146 561134
rect 231382 560898 240146 561134
rect 240382 560898 249146 561134
rect 249382 560898 258146 561134
rect 258382 560898 267146 561134
rect 267382 560898 269708 561134
rect 269944 560898 270360 561134
rect 270596 560898 271166 561134
rect 271402 560898 280166 561134
rect 280402 560898 289166 561134
rect 289402 560898 298166 561134
rect 298402 560898 307166 561134
rect 307402 560898 309728 561134
rect 309964 560898 311380 561134
rect 311616 560898 312186 561134
rect 312422 560898 321186 561134
rect 321422 560898 330186 561134
rect 330422 560898 339186 561134
rect 339422 560898 348186 561134
rect 348422 560898 350748 561134
rect 350984 560898 352400 561134
rect 352636 560898 353206 561134
rect 353442 560898 362206 561134
rect 362442 560898 371206 561134
rect 371442 560898 380206 561134
rect 380442 560898 389206 561134
rect 389442 560898 391768 561134
rect 392004 560898 392420 561134
rect 392656 560898 393226 561134
rect 393462 560898 402226 561134
rect 402462 560898 411226 561134
rect 411462 560898 420226 561134
rect 420462 560898 429226 561134
rect 429462 560898 431788 561134
rect 432024 560898 432440 561134
rect 432676 560898 433246 561134
rect 433482 560898 439792 561134
rect 440028 560898 457010 561134
rect 457246 560898 476652 561134
rect 476888 560898 571716 561134
rect 571952 560898 579470 561134
rect 579706 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 5382 543454
rect 5618 543218 127458 543454
rect 127694 543218 140656 543454
rect 140892 543218 141502 543454
rect 141738 543218 147288 543454
rect 147524 543218 149660 543454
rect 149896 543218 150506 543454
rect 150742 543218 159506 543454
rect 159742 543218 168506 543454
rect 168742 543218 177506 543454
rect 177742 543218 186506 543454
rect 186742 543218 188308 543454
rect 188544 543218 190680 543454
rect 190916 543218 191526 543454
rect 191762 543218 200526 543454
rect 200762 543218 209526 543454
rect 209762 543218 218526 543454
rect 218762 543218 227526 543454
rect 227762 543218 229328 543454
rect 229564 543218 230700 543454
rect 230936 543218 231546 543454
rect 231782 543218 240546 543454
rect 240782 543218 249546 543454
rect 249782 543218 258546 543454
rect 258782 543218 267546 543454
rect 267782 543218 269348 543454
rect 269584 543218 270720 543454
rect 270956 543218 271566 543454
rect 271802 543218 280566 543454
rect 280802 543218 289566 543454
rect 289802 543218 298566 543454
rect 298802 543218 307566 543454
rect 307802 543218 309368 543454
rect 309604 543218 311740 543454
rect 311976 543218 312586 543454
rect 312822 543218 321586 543454
rect 321822 543218 330586 543454
rect 330822 543218 339586 543454
rect 339822 543218 348586 543454
rect 348822 543218 350388 543454
rect 350624 543218 352760 543454
rect 352996 543218 353606 543454
rect 353842 543218 362606 543454
rect 362842 543218 371606 543454
rect 371842 543218 380606 543454
rect 380842 543218 389606 543454
rect 389842 543218 391408 543454
rect 391644 543218 392780 543454
rect 393016 543218 393626 543454
rect 393862 543218 402626 543454
rect 402862 543218 411626 543454
rect 411862 543218 420626 543454
rect 420862 543218 429626 543454
rect 429862 543218 431428 543454
rect 431664 543218 432800 543454
rect 433036 543218 433646 543454
rect 433882 543218 439432 543454
rect 439668 543218 456610 543454
rect 456846 543218 578670 543454
rect 578906 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 5382 543134
rect 5618 542898 127458 543134
rect 127694 542898 140656 543134
rect 140892 542898 141502 543134
rect 141738 542898 147288 543134
rect 147524 542898 149660 543134
rect 149896 542898 150506 543134
rect 150742 542898 159506 543134
rect 159742 542898 168506 543134
rect 168742 542898 177506 543134
rect 177742 542898 186506 543134
rect 186742 542898 188308 543134
rect 188544 542898 190680 543134
rect 190916 542898 191526 543134
rect 191762 542898 200526 543134
rect 200762 542898 209526 543134
rect 209762 542898 218526 543134
rect 218762 542898 227526 543134
rect 227762 542898 229328 543134
rect 229564 542898 230700 543134
rect 230936 542898 231546 543134
rect 231782 542898 240546 543134
rect 240782 542898 249546 543134
rect 249782 542898 258546 543134
rect 258782 542898 267546 543134
rect 267782 542898 269348 543134
rect 269584 542898 270720 543134
rect 270956 542898 271566 543134
rect 271802 542898 280566 543134
rect 280802 542898 289566 543134
rect 289802 542898 298566 543134
rect 298802 542898 307566 543134
rect 307802 542898 309368 543134
rect 309604 542898 311740 543134
rect 311976 542898 312586 543134
rect 312822 542898 321586 543134
rect 321822 542898 330586 543134
rect 330822 542898 339586 543134
rect 339822 542898 348586 543134
rect 348822 542898 350388 543134
rect 350624 542898 352760 543134
rect 352996 542898 353606 543134
rect 353842 542898 362606 543134
rect 362842 542898 371606 543134
rect 371842 542898 380606 543134
rect 380842 542898 389606 543134
rect 389842 542898 391408 543134
rect 391644 542898 392780 543134
rect 393016 542898 393626 543134
rect 393862 542898 402626 543134
rect 402862 542898 411626 543134
rect 411862 542898 420626 543134
rect 420862 542898 429626 543134
rect 429862 542898 431428 543134
rect 431664 542898 432800 543134
rect 433036 542898 433646 543134
rect 433882 542898 439432 543134
rect 439668 542898 456610 543134
rect 456846 542898 578670 543134
rect 578906 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 4582 525454
rect 4818 525218 127058 525454
rect 127294 525218 140296 525454
rect 140532 525218 141102 525454
rect 141338 525218 147648 525454
rect 147884 525218 149300 525454
rect 149536 525218 150106 525454
rect 150342 525218 159106 525454
rect 159342 525218 168106 525454
rect 168342 525218 177106 525454
rect 177342 525218 186106 525454
rect 186342 525218 188668 525454
rect 188904 525218 190320 525454
rect 190556 525218 191126 525454
rect 191362 525218 200126 525454
rect 200362 525218 209126 525454
rect 209362 525218 218126 525454
rect 218362 525218 227126 525454
rect 227362 525218 229688 525454
rect 229924 525218 230340 525454
rect 230576 525218 231146 525454
rect 231382 525218 240146 525454
rect 240382 525218 249146 525454
rect 249382 525218 258146 525454
rect 258382 525218 267146 525454
rect 267382 525218 269708 525454
rect 269944 525218 270360 525454
rect 270596 525218 271166 525454
rect 271402 525218 280166 525454
rect 280402 525218 289166 525454
rect 289402 525218 298166 525454
rect 298402 525218 307166 525454
rect 307402 525218 309728 525454
rect 309964 525218 311380 525454
rect 311616 525218 312186 525454
rect 312422 525218 321186 525454
rect 321422 525218 330186 525454
rect 330422 525218 339186 525454
rect 339422 525218 348186 525454
rect 348422 525218 350748 525454
rect 350984 525218 352400 525454
rect 352636 525218 353206 525454
rect 353442 525218 362206 525454
rect 362442 525218 371206 525454
rect 371442 525218 380206 525454
rect 380442 525218 389206 525454
rect 389442 525218 391768 525454
rect 392004 525218 392420 525454
rect 392656 525218 393226 525454
rect 393462 525218 402226 525454
rect 402462 525218 411226 525454
rect 411462 525218 420226 525454
rect 420462 525218 429226 525454
rect 429462 525218 431788 525454
rect 432024 525218 432440 525454
rect 432676 525218 433246 525454
rect 433482 525218 439792 525454
rect 440028 525218 457010 525454
rect 457246 525218 579470 525454
rect 579706 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 4582 525134
rect 4818 524898 127058 525134
rect 127294 524898 140296 525134
rect 140532 524898 141102 525134
rect 141338 524898 147648 525134
rect 147884 524898 149300 525134
rect 149536 524898 150106 525134
rect 150342 524898 159106 525134
rect 159342 524898 168106 525134
rect 168342 524898 177106 525134
rect 177342 524898 186106 525134
rect 186342 524898 188668 525134
rect 188904 524898 190320 525134
rect 190556 524898 191126 525134
rect 191362 524898 200126 525134
rect 200362 524898 209126 525134
rect 209362 524898 218126 525134
rect 218362 524898 227126 525134
rect 227362 524898 229688 525134
rect 229924 524898 230340 525134
rect 230576 524898 231146 525134
rect 231382 524898 240146 525134
rect 240382 524898 249146 525134
rect 249382 524898 258146 525134
rect 258382 524898 267146 525134
rect 267382 524898 269708 525134
rect 269944 524898 270360 525134
rect 270596 524898 271166 525134
rect 271402 524898 280166 525134
rect 280402 524898 289166 525134
rect 289402 524898 298166 525134
rect 298402 524898 307166 525134
rect 307402 524898 309728 525134
rect 309964 524898 311380 525134
rect 311616 524898 312186 525134
rect 312422 524898 321186 525134
rect 321422 524898 330186 525134
rect 330422 524898 339186 525134
rect 339422 524898 348186 525134
rect 348422 524898 350748 525134
rect 350984 524898 352400 525134
rect 352636 524898 353206 525134
rect 353442 524898 362206 525134
rect 362442 524898 371206 525134
rect 371442 524898 380206 525134
rect 380442 524898 389206 525134
rect 389442 524898 391768 525134
rect 392004 524898 392420 525134
rect 392656 524898 393226 525134
rect 393462 524898 402226 525134
rect 402462 524898 411226 525134
rect 411462 524898 420226 525134
rect 420462 524898 429226 525134
rect 429462 524898 431788 525134
rect 432024 524898 432440 525134
rect 432676 524898 433246 525134
rect 433482 524898 439792 525134
rect 440028 524898 457010 525134
rect 457246 524898 579470 525134
rect 579706 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 5382 507454
rect 5618 507218 127458 507454
rect 127694 507218 140656 507454
rect 140892 507218 141502 507454
rect 141738 507218 147288 507454
rect 147524 507218 149660 507454
rect 149896 507218 150506 507454
rect 150742 507218 159506 507454
rect 159742 507218 168506 507454
rect 168742 507218 177506 507454
rect 177742 507218 186506 507454
rect 186742 507218 188308 507454
rect 188544 507218 190680 507454
rect 190916 507218 191526 507454
rect 191762 507218 200526 507454
rect 200762 507218 209526 507454
rect 209762 507218 218526 507454
rect 218762 507218 227526 507454
rect 227762 507218 229328 507454
rect 229564 507218 230700 507454
rect 230936 507218 231546 507454
rect 231782 507218 240546 507454
rect 240782 507218 249546 507454
rect 249782 507218 258546 507454
rect 258782 507218 267546 507454
rect 267782 507218 269348 507454
rect 269584 507218 270720 507454
rect 270956 507218 271566 507454
rect 271802 507218 280566 507454
rect 280802 507218 289566 507454
rect 289802 507218 298566 507454
rect 298802 507218 307566 507454
rect 307802 507218 309368 507454
rect 309604 507218 311740 507454
rect 311976 507218 312586 507454
rect 312822 507218 321586 507454
rect 321822 507218 330586 507454
rect 330822 507218 339586 507454
rect 339822 507218 348586 507454
rect 348822 507218 350388 507454
rect 350624 507218 352760 507454
rect 352996 507218 353606 507454
rect 353842 507218 362606 507454
rect 362842 507218 371606 507454
rect 371842 507218 380606 507454
rect 380842 507218 389606 507454
rect 389842 507218 391408 507454
rect 391644 507218 392780 507454
rect 393016 507218 393626 507454
rect 393862 507218 402626 507454
rect 402862 507218 411626 507454
rect 411862 507218 420626 507454
rect 420862 507218 429626 507454
rect 429862 507218 431428 507454
rect 431664 507218 432800 507454
rect 433036 507218 433646 507454
rect 433882 507218 439432 507454
rect 439668 507218 456610 507454
rect 456846 507218 578670 507454
rect 578906 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 5382 507134
rect 5618 506898 127458 507134
rect 127694 506898 140656 507134
rect 140892 506898 141502 507134
rect 141738 506898 147288 507134
rect 147524 506898 149660 507134
rect 149896 506898 150506 507134
rect 150742 506898 159506 507134
rect 159742 506898 168506 507134
rect 168742 506898 177506 507134
rect 177742 506898 186506 507134
rect 186742 506898 188308 507134
rect 188544 506898 190680 507134
rect 190916 506898 191526 507134
rect 191762 506898 200526 507134
rect 200762 506898 209526 507134
rect 209762 506898 218526 507134
rect 218762 506898 227526 507134
rect 227762 506898 229328 507134
rect 229564 506898 230700 507134
rect 230936 506898 231546 507134
rect 231782 506898 240546 507134
rect 240782 506898 249546 507134
rect 249782 506898 258546 507134
rect 258782 506898 267546 507134
rect 267782 506898 269348 507134
rect 269584 506898 270720 507134
rect 270956 506898 271566 507134
rect 271802 506898 280566 507134
rect 280802 506898 289566 507134
rect 289802 506898 298566 507134
rect 298802 506898 307566 507134
rect 307802 506898 309368 507134
rect 309604 506898 311740 507134
rect 311976 506898 312586 507134
rect 312822 506898 321586 507134
rect 321822 506898 330586 507134
rect 330822 506898 339586 507134
rect 339822 506898 348586 507134
rect 348822 506898 350388 507134
rect 350624 506898 352760 507134
rect 352996 506898 353606 507134
rect 353842 506898 362606 507134
rect 362842 506898 371606 507134
rect 371842 506898 380606 507134
rect 380842 506898 389606 507134
rect 389842 506898 391408 507134
rect 391644 506898 392780 507134
rect 393016 506898 393626 507134
rect 393862 506898 402626 507134
rect 402862 506898 411626 507134
rect 411862 506898 420626 507134
rect 420862 506898 429626 507134
rect 429862 506898 431428 507134
rect 431664 506898 432800 507134
rect 433036 506898 433646 507134
rect 433882 506898 439432 507134
rect 439668 506898 456610 507134
rect 456846 506898 578670 507134
rect 578906 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 4582 489454
rect 4818 489218 12618 489454
rect 12854 489218 14040 489454
rect 14276 489218 23040 489454
rect 23276 489218 32040 489454
rect 32276 489218 41040 489454
rect 41276 489218 50040 489454
rect 50276 489218 59040 489454
rect 59276 489218 68040 489454
rect 68276 489218 77040 489454
rect 77276 489218 86040 489454
rect 86276 489218 95040 489454
rect 95276 489218 104040 489454
rect 104276 489218 113040 489454
rect 113276 489218 121226 489454
rect 121462 489218 127058 489454
rect 127294 489218 140296 489454
rect 140532 489218 141102 489454
rect 141338 489218 147648 489454
rect 147884 489218 149300 489454
rect 149536 489218 150106 489454
rect 150342 489218 159106 489454
rect 159342 489218 168106 489454
rect 168342 489218 177106 489454
rect 177342 489218 186106 489454
rect 186342 489218 188668 489454
rect 188904 489218 189768 489454
rect 190004 489218 190320 489454
rect 190556 489218 191126 489454
rect 191362 489218 200126 489454
rect 200362 489218 209126 489454
rect 209362 489218 218126 489454
rect 218362 489218 227126 489454
rect 227362 489218 229688 489454
rect 229924 489218 230340 489454
rect 230576 489218 231146 489454
rect 231382 489218 240146 489454
rect 240382 489218 249146 489454
rect 249382 489218 258146 489454
rect 258382 489218 267146 489454
rect 267382 489218 269708 489454
rect 269944 489218 270360 489454
rect 270596 489218 271166 489454
rect 271402 489218 280166 489454
rect 280402 489218 289166 489454
rect 289402 489218 298166 489454
rect 298402 489218 307166 489454
rect 307402 489218 309728 489454
rect 309964 489218 311380 489454
rect 311616 489218 312186 489454
rect 312422 489218 321186 489454
rect 321422 489218 330186 489454
rect 330422 489218 339186 489454
rect 339422 489218 348186 489454
rect 348422 489218 350748 489454
rect 350984 489218 352400 489454
rect 352636 489218 353206 489454
rect 353442 489218 362206 489454
rect 362442 489218 371206 489454
rect 371442 489218 380206 489454
rect 380442 489218 389206 489454
rect 389442 489218 391768 489454
rect 392004 489218 392420 489454
rect 392656 489218 393226 489454
rect 393462 489218 402226 489454
rect 402462 489218 411226 489454
rect 411462 489218 420226 489454
rect 420462 489218 429226 489454
rect 429462 489218 431788 489454
rect 432024 489218 432440 489454
rect 432676 489218 433246 489454
rect 433482 489218 439792 489454
rect 440028 489218 457010 489454
rect 457246 489218 462842 489454
rect 463078 489218 471028 489454
rect 471264 489218 480028 489454
rect 480264 489218 489028 489454
rect 489264 489218 498028 489454
rect 498264 489218 507028 489454
rect 507264 489218 516028 489454
rect 516264 489218 525028 489454
rect 525264 489218 534028 489454
rect 534264 489218 543028 489454
rect 543264 489218 552028 489454
rect 552264 489218 561028 489454
rect 561264 489218 570028 489454
rect 570264 489218 571450 489454
rect 571686 489218 579470 489454
rect 579706 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 4582 489134
rect 4818 488898 12618 489134
rect 12854 488898 14040 489134
rect 14276 488898 23040 489134
rect 23276 488898 32040 489134
rect 32276 488898 41040 489134
rect 41276 488898 50040 489134
rect 50276 488898 59040 489134
rect 59276 488898 68040 489134
rect 68276 488898 77040 489134
rect 77276 488898 86040 489134
rect 86276 488898 95040 489134
rect 95276 488898 104040 489134
rect 104276 488898 113040 489134
rect 113276 488898 121226 489134
rect 121462 488898 127058 489134
rect 127294 488898 140296 489134
rect 140532 488898 141102 489134
rect 141338 488898 147648 489134
rect 147884 488898 149300 489134
rect 149536 488898 150106 489134
rect 150342 488898 159106 489134
rect 159342 488898 168106 489134
rect 168342 488898 177106 489134
rect 177342 488898 186106 489134
rect 186342 488898 188668 489134
rect 188904 488898 189768 489134
rect 190004 488898 190320 489134
rect 190556 488898 191126 489134
rect 191362 488898 200126 489134
rect 200362 488898 209126 489134
rect 209362 488898 218126 489134
rect 218362 488898 227126 489134
rect 227362 488898 229688 489134
rect 229924 488898 230340 489134
rect 230576 488898 231146 489134
rect 231382 488898 240146 489134
rect 240382 488898 249146 489134
rect 249382 488898 258146 489134
rect 258382 488898 267146 489134
rect 267382 488898 269708 489134
rect 269944 488898 270360 489134
rect 270596 488898 271166 489134
rect 271402 488898 280166 489134
rect 280402 488898 289166 489134
rect 289402 488898 298166 489134
rect 298402 488898 307166 489134
rect 307402 488898 309728 489134
rect 309964 488898 311380 489134
rect 311616 488898 312186 489134
rect 312422 488898 321186 489134
rect 321422 488898 330186 489134
rect 330422 488898 339186 489134
rect 339422 488898 348186 489134
rect 348422 488898 350748 489134
rect 350984 488898 352400 489134
rect 352636 488898 353206 489134
rect 353442 488898 362206 489134
rect 362442 488898 371206 489134
rect 371442 488898 380206 489134
rect 380442 488898 389206 489134
rect 389442 488898 391768 489134
rect 392004 488898 392420 489134
rect 392656 488898 393226 489134
rect 393462 488898 402226 489134
rect 402462 488898 411226 489134
rect 411462 488898 420226 489134
rect 420462 488898 429226 489134
rect 429462 488898 431788 489134
rect 432024 488898 432440 489134
rect 432676 488898 433246 489134
rect 433482 488898 439792 489134
rect 440028 488898 457010 489134
rect 457246 488898 462842 489134
rect 463078 488898 471028 489134
rect 471264 488898 480028 489134
rect 480264 488898 489028 489134
rect 489264 488898 498028 489134
rect 498264 488898 507028 489134
rect 507264 488898 516028 489134
rect 516264 488898 525028 489134
rect 525264 488898 534028 489134
rect 534264 488898 543028 489134
rect 543264 488898 552028 489134
rect 552264 488898 561028 489134
rect 561264 488898 570028 489134
rect 570264 488898 571450 489134
rect 571686 488898 579470 489134
rect 579706 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 5382 471454
rect 5618 471218 13218 471454
rect 13454 471218 14420 471454
rect 14656 471218 23420 471454
rect 23656 471218 32420 471454
rect 32656 471218 41420 471454
rect 41656 471218 50420 471454
rect 50656 471218 59420 471454
rect 59656 471218 68420 471454
rect 68656 471218 77420 471454
rect 77656 471218 86420 471454
rect 86656 471218 95420 471454
rect 95656 471218 104420 471454
rect 104656 471218 113420 471454
rect 113656 471218 120626 471454
rect 120862 471218 127458 471454
rect 127694 471218 140656 471454
rect 140892 471218 141502 471454
rect 141738 471218 147288 471454
rect 147524 471218 149660 471454
rect 149896 471218 150506 471454
rect 150742 471218 159506 471454
rect 159742 471218 168506 471454
rect 168742 471218 177506 471454
rect 177742 471218 186506 471454
rect 186742 471218 188308 471454
rect 188544 471218 190680 471454
rect 190916 471218 191526 471454
rect 191762 471218 200526 471454
rect 200762 471218 209526 471454
rect 209762 471218 218526 471454
rect 218762 471218 227526 471454
rect 227762 471218 229328 471454
rect 229564 471218 230700 471454
rect 230936 471218 231546 471454
rect 231782 471218 240546 471454
rect 240782 471218 249546 471454
rect 249782 471218 258546 471454
rect 258782 471218 267546 471454
rect 267782 471218 269348 471454
rect 269584 471218 270720 471454
rect 270956 471218 271566 471454
rect 271802 471218 280566 471454
rect 280802 471218 289566 471454
rect 289802 471218 298566 471454
rect 298802 471218 307566 471454
rect 307802 471218 309368 471454
rect 309604 471218 311740 471454
rect 311976 471218 312586 471454
rect 312822 471218 321586 471454
rect 321822 471218 330586 471454
rect 330822 471218 339586 471454
rect 339822 471218 348586 471454
rect 348822 471218 350388 471454
rect 350624 471218 352760 471454
rect 352996 471218 353606 471454
rect 353842 471218 362606 471454
rect 362842 471218 371606 471454
rect 371842 471218 380606 471454
rect 380842 471218 389606 471454
rect 389842 471218 391408 471454
rect 391644 471218 392780 471454
rect 393016 471218 393626 471454
rect 393862 471218 402626 471454
rect 402862 471218 411626 471454
rect 411862 471218 420626 471454
rect 420862 471218 429626 471454
rect 429862 471218 431428 471454
rect 431664 471218 432800 471454
rect 433036 471218 433646 471454
rect 433882 471218 439432 471454
rect 439668 471218 456610 471454
rect 456846 471218 463442 471454
rect 463678 471218 470648 471454
rect 470884 471218 479648 471454
rect 479884 471218 488648 471454
rect 488884 471218 497648 471454
rect 497884 471218 506648 471454
rect 506884 471218 515648 471454
rect 515884 471218 524648 471454
rect 524884 471218 533648 471454
rect 533884 471218 542648 471454
rect 542884 471218 551648 471454
rect 551884 471218 560648 471454
rect 560884 471218 569648 471454
rect 569884 471218 570850 471454
rect 571086 471218 578670 471454
rect 578906 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 5382 471134
rect 5618 470898 13218 471134
rect 13454 470898 14420 471134
rect 14656 470898 23420 471134
rect 23656 470898 32420 471134
rect 32656 470898 41420 471134
rect 41656 470898 50420 471134
rect 50656 470898 59420 471134
rect 59656 470898 68420 471134
rect 68656 470898 77420 471134
rect 77656 470898 86420 471134
rect 86656 470898 95420 471134
rect 95656 470898 104420 471134
rect 104656 470898 113420 471134
rect 113656 470898 120626 471134
rect 120862 470898 127458 471134
rect 127694 470898 140656 471134
rect 140892 470898 141502 471134
rect 141738 470898 147288 471134
rect 147524 470898 149660 471134
rect 149896 470898 150506 471134
rect 150742 470898 159506 471134
rect 159742 470898 168506 471134
rect 168742 470898 177506 471134
rect 177742 470898 186506 471134
rect 186742 470898 188308 471134
rect 188544 470898 190680 471134
rect 190916 470898 191526 471134
rect 191762 470898 200526 471134
rect 200762 470898 209526 471134
rect 209762 470898 218526 471134
rect 218762 470898 227526 471134
rect 227762 470898 229328 471134
rect 229564 470898 230700 471134
rect 230936 470898 231546 471134
rect 231782 470898 240546 471134
rect 240782 470898 249546 471134
rect 249782 470898 258546 471134
rect 258782 470898 267546 471134
rect 267782 470898 269348 471134
rect 269584 470898 270720 471134
rect 270956 470898 271566 471134
rect 271802 470898 280566 471134
rect 280802 470898 289566 471134
rect 289802 470898 298566 471134
rect 298802 470898 307566 471134
rect 307802 470898 309368 471134
rect 309604 470898 311740 471134
rect 311976 470898 312586 471134
rect 312822 470898 321586 471134
rect 321822 470898 330586 471134
rect 330822 470898 339586 471134
rect 339822 470898 348586 471134
rect 348822 470898 350388 471134
rect 350624 470898 352760 471134
rect 352996 470898 353606 471134
rect 353842 470898 362606 471134
rect 362842 470898 371606 471134
rect 371842 470898 380606 471134
rect 380842 470898 389606 471134
rect 389842 470898 391408 471134
rect 391644 470898 392780 471134
rect 393016 470898 393626 471134
rect 393862 470898 402626 471134
rect 402862 470898 411626 471134
rect 411862 470898 420626 471134
rect 420862 470898 429626 471134
rect 429862 470898 431428 471134
rect 431664 470898 432800 471134
rect 433036 470898 433646 471134
rect 433882 470898 439432 471134
rect 439668 470898 456610 471134
rect 456846 470898 463442 471134
rect 463678 470898 470648 471134
rect 470884 470898 479648 471134
rect 479884 470898 488648 471134
rect 488884 470898 497648 471134
rect 497884 470898 506648 471134
rect 506884 470898 515648 471134
rect 515884 470898 524648 471134
rect 524884 470898 533648 471134
rect 533884 470898 542648 471134
rect 542884 470898 551648 471134
rect 551884 470898 560648 471134
rect 560884 470898 569648 471134
rect 569884 470898 570850 471134
rect 571086 470898 578670 471134
rect 578906 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 4582 453454
rect 4818 453218 12618 453454
rect 12854 453218 14040 453454
rect 14276 453218 23040 453454
rect 23276 453218 32040 453454
rect 32276 453218 41040 453454
rect 41276 453218 50040 453454
rect 50276 453218 59040 453454
rect 59276 453218 68040 453454
rect 68276 453218 77040 453454
rect 77276 453218 86040 453454
rect 86276 453218 95040 453454
rect 95276 453218 104040 453454
rect 104276 453218 113040 453454
rect 113276 453218 121226 453454
rect 121462 453218 127058 453454
rect 127294 453218 140296 453454
rect 140532 453218 141102 453454
rect 141338 453218 147648 453454
rect 147884 453218 149300 453454
rect 149536 453218 150106 453454
rect 150342 453218 159106 453454
rect 159342 453218 168106 453454
rect 168342 453218 177106 453454
rect 177342 453218 186106 453454
rect 186342 453218 188668 453454
rect 188904 453218 190320 453454
rect 190556 453218 191126 453454
rect 191362 453218 200126 453454
rect 200362 453218 209126 453454
rect 209362 453218 218126 453454
rect 218362 453218 227126 453454
rect 227362 453218 229688 453454
rect 229924 453218 230340 453454
rect 230576 453218 231146 453454
rect 231382 453218 240146 453454
rect 240382 453218 249146 453454
rect 249382 453218 258146 453454
rect 258382 453218 267146 453454
rect 267382 453218 269708 453454
rect 269944 453218 270360 453454
rect 270596 453218 271166 453454
rect 271402 453218 280166 453454
rect 280402 453218 289166 453454
rect 289402 453218 298166 453454
rect 298402 453218 307166 453454
rect 307402 453218 309728 453454
rect 309964 453218 311380 453454
rect 311616 453218 312186 453454
rect 312422 453218 321186 453454
rect 321422 453218 330186 453454
rect 330422 453218 339186 453454
rect 339422 453218 348186 453454
rect 348422 453218 350748 453454
rect 350984 453218 352400 453454
rect 352636 453218 353206 453454
rect 353442 453218 362206 453454
rect 362442 453218 371206 453454
rect 371442 453218 380206 453454
rect 380442 453218 389206 453454
rect 389442 453218 391768 453454
rect 392004 453218 392420 453454
rect 392656 453218 393226 453454
rect 393462 453218 402226 453454
rect 402462 453218 411226 453454
rect 411462 453218 420226 453454
rect 420462 453218 429226 453454
rect 429462 453218 431788 453454
rect 432024 453218 432440 453454
rect 432676 453218 433246 453454
rect 433482 453218 439792 453454
rect 440028 453218 457010 453454
rect 457246 453218 462842 453454
rect 463078 453218 471028 453454
rect 471264 453218 480028 453454
rect 480264 453218 489028 453454
rect 489264 453218 498028 453454
rect 498264 453218 507028 453454
rect 507264 453218 516028 453454
rect 516264 453218 525028 453454
rect 525264 453218 534028 453454
rect 534264 453218 543028 453454
rect 543264 453218 552028 453454
rect 552264 453218 561028 453454
rect 561264 453218 570028 453454
rect 570264 453218 571450 453454
rect 571686 453218 579470 453454
rect 579706 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 4582 453134
rect 4818 452898 12618 453134
rect 12854 452898 14040 453134
rect 14276 452898 23040 453134
rect 23276 452898 32040 453134
rect 32276 452898 41040 453134
rect 41276 452898 50040 453134
rect 50276 452898 59040 453134
rect 59276 452898 68040 453134
rect 68276 452898 77040 453134
rect 77276 452898 86040 453134
rect 86276 452898 95040 453134
rect 95276 452898 104040 453134
rect 104276 452898 113040 453134
rect 113276 452898 121226 453134
rect 121462 452898 127058 453134
rect 127294 452898 140296 453134
rect 140532 452898 141102 453134
rect 141338 452898 147648 453134
rect 147884 452898 149300 453134
rect 149536 452898 150106 453134
rect 150342 452898 159106 453134
rect 159342 452898 168106 453134
rect 168342 452898 177106 453134
rect 177342 452898 186106 453134
rect 186342 452898 188668 453134
rect 188904 452898 190320 453134
rect 190556 452898 191126 453134
rect 191362 452898 200126 453134
rect 200362 452898 209126 453134
rect 209362 452898 218126 453134
rect 218362 452898 227126 453134
rect 227362 452898 229688 453134
rect 229924 452898 230340 453134
rect 230576 452898 231146 453134
rect 231382 452898 240146 453134
rect 240382 452898 249146 453134
rect 249382 452898 258146 453134
rect 258382 452898 267146 453134
rect 267382 452898 269708 453134
rect 269944 452898 270360 453134
rect 270596 452898 271166 453134
rect 271402 452898 280166 453134
rect 280402 452898 289166 453134
rect 289402 452898 298166 453134
rect 298402 452898 307166 453134
rect 307402 452898 309728 453134
rect 309964 452898 311380 453134
rect 311616 452898 312186 453134
rect 312422 452898 321186 453134
rect 321422 452898 330186 453134
rect 330422 452898 339186 453134
rect 339422 452898 348186 453134
rect 348422 452898 350748 453134
rect 350984 452898 352400 453134
rect 352636 452898 353206 453134
rect 353442 452898 362206 453134
rect 362442 452898 371206 453134
rect 371442 452898 380206 453134
rect 380442 452898 389206 453134
rect 389442 452898 391768 453134
rect 392004 452898 392420 453134
rect 392656 452898 393226 453134
rect 393462 452898 402226 453134
rect 402462 452898 411226 453134
rect 411462 452898 420226 453134
rect 420462 452898 429226 453134
rect 429462 452898 431788 453134
rect 432024 452898 432440 453134
rect 432676 452898 433246 453134
rect 433482 452898 439792 453134
rect 440028 452898 457010 453134
rect 457246 452898 462842 453134
rect 463078 452898 471028 453134
rect 471264 452898 480028 453134
rect 480264 452898 489028 453134
rect 489264 452898 498028 453134
rect 498264 452898 507028 453134
rect 507264 452898 516028 453134
rect 516264 452898 525028 453134
rect 525264 452898 534028 453134
rect 534264 452898 543028 453134
rect 543264 452898 552028 453134
rect 552264 452898 561028 453134
rect 561264 452898 570028 453134
rect 570264 452898 571450 453134
rect 571686 452898 579470 453134
rect 579706 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 5382 435454
rect 5618 435218 13218 435454
rect 13454 435218 14420 435454
rect 14656 435218 23420 435454
rect 23656 435218 32420 435454
rect 32656 435218 41420 435454
rect 41656 435218 50420 435454
rect 50656 435218 59420 435454
rect 59656 435218 68420 435454
rect 68656 435218 77420 435454
rect 77656 435218 86420 435454
rect 86656 435218 95420 435454
rect 95656 435218 104420 435454
rect 104656 435218 113420 435454
rect 113656 435218 120626 435454
rect 120862 435218 127458 435454
rect 127694 435218 140656 435454
rect 140892 435218 147288 435454
rect 147524 435218 149660 435454
rect 149896 435218 150506 435454
rect 150742 435218 159506 435454
rect 159742 435218 168506 435454
rect 168742 435218 177506 435454
rect 177742 435218 186506 435454
rect 186742 435218 188308 435454
rect 188544 435218 190680 435454
rect 190916 435218 229328 435454
rect 229564 435218 230700 435454
rect 230936 435218 269348 435454
rect 269584 435218 270720 435454
rect 270956 435218 309368 435454
rect 309604 435218 311740 435454
rect 311976 435218 312586 435454
rect 312822 435218 321586 435454
rect 321822 435218 330586 435454
rect 330822 435218 339586 435454
rect 339822 435218 348586 435454
rect 348822 435218 350388 435454
rect 350624 435218 352760 435454
rect 352996 435218 391408 435454
rect 391644 435218 392780 435454
rect 393016 435218 431428 435454
rect 431664 435218 432800 435454
rect 433036 435218 439432 435454
rect 439668 435218 456610 435454
rect 456846 435218 463442 435454
rect 463678 435218 470648 435454
rect 470884 435218 479648 435454
rect 479884 435218 488648 435454
rect 488884 435218 497648 435454
rect 497884 435218 506648 435454
rect 506884 435218 515648 435454
rect 515884 435218 524648 435454
rect 524884 435218 533648 435454
rect 533884 435218 542648 435454
rect 542884 435218 551648 435454
rect 551884 435218 560648 435454
rect 560884 435218 569648 435454
rect 569884 435218 570850 435454
rect 571086 435218 578670 435454
rect 578906 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 5382 435134
rect 5618 434898 13218 435134
rect 13454 434898 14420 435134
rect 14656 434898 23420 435134
rect 23656 434898 32420 435134
rect 32656 434898 41420 435134
rect 41656 434898 50420 435134
rect 50656 434898 59420 435134
rect 59656 434898 68420 435134
rect 68656 434898 77420 435134
rect 77656 434898 86420 435134
rect 86656 434898 95420 435134
rect 95656 434898 104420 435134
rect 104656 434898 113420 435134
rect 113656 434898 120626 435134
rect 120862 434898 127458 435134
rect 127694 434898 140656 435134
rect 140892 434898 147288 435134
rect 147524 434898 149660 435134
rect 149896 434898 150506 435134
rect 150742 434898 159506 435134
rect 159742 434898 168506 435134
rect 168742 434898 177506 435134
rect 177742 434898 186506 435134
rect 186742 434898 188308 435134
rect 188544 434898 190680 435134
rect 190916 434898 229328 435134
rect 229564 434898 230700 435134
rect 230936 434898 269348 435134
rect 269584 434898 270720 435134
rect 270956 434898 309368 435134
rect 309604 434898 311740 435134
rect 311976 434898 312586 435134
rect 312822 434898 321586 435134
rect 321822 434898 330586 435134
rect 330822 434898 339586 435134
rect 339822 434898 348586 435134
rect 348822 434898 350388 435134
rect 350624 434898 352760 435134
rect 352996 434898 391408 435134
rect 391644 434898 392780 435134
rect 393016 434898 431428 435134
rect 431664 434898 432800 435134
rect 433036 434898 439432 435134
rect 439668 434898 456610 435134
rect 456846 434898 463442 435134
rect 463678 434898 470648 435134
rect 470884 434898 479648 435134
rect 479884 434898 488648 435134
rect 488884 434898 497648 435134
rect 497884 434898 506648 435134
rect 506884 434898 515648 435134
rect 515884 434898 524648 435134
rect 524884 434898 533648 435134
rect 533884 434898 542648 435134
rect 542884 434898 551648 435134
rect 551884 434898 560648 435134
rect 560884 434898 569648 435134
rect 569884 434898 570850 435134
rect 571086 434898 578670 435134
rect 578906 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 4582 417454
rect 4818 417218 12618 417454
rect 12854 417218 14040 417454
rect 14276 417218 23040 417454
rect 23276 417218 32040 417454
rect 32276 417218 41040 417454
rect 41276 417218 50040 417454
rect 50276 417218 59040 417454
rect 59276 417218 68040 417454
rect 68276 417218 77040 417454
rect 77276 417218 86040 417454
rect 86276 417218 95040 417454
rect 95276 417218 104040 417454
rect 104276 417218 113040 417454
rect 113276 417218 121226 417454
rect 121462 417218 127058 417454
rect 127294 417218 140296 417454
rect 140532 417218 141102 417454
rect 141338 417218 147648 417454
rect 147884 417218 149300 417454
rect 149536 417218 150106 417454
rect 150342 417218 159106 417454
rect 159342 417218 168106 417454
rect 168342 417218 177106 417454
rect 177342 417218 186106 417454
rect 186342 417218 188668 417454
rect 188904 417218 189768 417454
rect 190004 417218 190320 417454
rect 190556 417218 191126 417454
rect 191362 417218 200126 417454
rect 200362 417218 209126 417454
rect 209362 417218 218126 417454
rect 218362 417218 227126 417454
rect 227362 417218 229688 417454
rect 229924 417218 230340 417454
rect 230576 417218 231146 417454
rect 231382 417218 240146 417454
rect 240382 417218 249146 417454
rect 249382 417218 258146 417454
rect 258382 417218 267146 417454
rect 267382 417218 269708 417454
rect 269944 417218 270360 417454
rect 270596 417218 271166 417454
rect 271402 417218 280166 417454
rect 280402 417218 289166 417454
rect 289402 417218 298166 417454
rect 298402 417218 307166 417454
rect 307402 417218 309728 417454
rect 309964 417218 311380 417454
rect 311616 417218 312186 417454
rect 312422 417218 321186 417454
rect 321422 417218 330186 417454
rect 330422 417218 339186 417454
rect 339422 417218 348186 417454
rect 348422 417218 350748 417454
rect 350984 417218 352400 417454
rect 352636 417218 353206 417454
rect 353442 417218 362206 417454
rect 362442 417218 371206 417454
rect 371442 417218 380206 417454
rect 380442 417218 389206 417454
rect 389442 417218 391768 417454
rect 392004 417218 392420 417454
rect 392656 417218 393226 417454
rect 393462 417218 402226 417454
rect 402462 417218 411226 417454
rect 411462 417218 420226 417454
rect 420462 417218 429226 417454
rect 429462 417218 431788 417454
rect 432024 417218 432440 417454
rect 432676 417218 433246 417454
rect 433482 417218 439792 417454
rect 440028 417218 457010 417454
rect 457246 417218 462842 417454
rect 463078 417218 471028 417454
rect 471264 417218 480028 417454
rect 480264 417218 489028 417454
rect 489264 417218 498028 417454
rect 498264 417218 507028 417454
rect 507264 417218 516028 417454
rect 516264 417218 525028 417454
rect 525264 417218 534028 417454
rect 534264 417218 543028 417454
rect 543264 417218 552028 417454
rect 552264 417218 561028 417454
rect 561264 417218 570028 417454
rect 570264 417218 571450 417454
rect 571686 417218 579470 417454
rect 579706 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 4582 417134
rect 4818 416898 12618 417134
rect 12854 416898 14040 417134
rect 14276 416898 23040 417134
rect 23276 416898 32040 417134
rect 32276 416898 41040 417134
rect 41276 416898 50040 417134
rect 50276 416898 59040 417134
rect 59276 416898 68040 417134
rect 68276 416898 77040 417134
rect 77276 416898 86040 417134
rect 86276 416898 95040 417134
rect 95276 416898 104040 417134
rect 104276 416898 113040 417134
rect 113276 416898 121226 417134
rect 121462 416898 127058 417134
rect 127294 416898 140296 417134
rect 140532 416898 141102 417134
rect 141338 416898 147648 417134
rect 147884 416898 149300 417134
rect 149536 416898 150106 417134
rect 150342 416898 159106 417134
rect 159342 416898 168106 417134
rect 168342 416898 177106 417134
rect 177342 416898 186106 417134
rect 186342 416898 188668 417134
rect 188904 416898 189768 417134
rect 190004 416898 190320 417134
rect 190556 416898 191126 417134
rect 191362 416898 200126 417134
rect 200362 416898 209126 417134
rect 209362 416898 218126 417134
rect 218362 416898 227126 417134
rect 227362 416898 229688 417134
rect 229924 416898 230340 417134
rect 230576 416898 231146 417134
rect 231382 416898 240146 417134
rect 240382 416898 249146 417134
rect 249382 416898 258146 417134
rect 258382 416898 267146 417134
rect 267382 416898 269708 417134
rect 269944 416898 270360 417134
rect 270596 416898 271166 417134
rect 271402 416898 280166 417134
rect 280402 416898 289166 417134
rect 289402 416898 298166 417134
rect 298402 416898 307166 417134
rect 307402 416898 309728 417134
rect 309964 416898 311380 417134
rect 311616 416898 312186 417134
rect 312422 416898 321186 417134
rect 321422 416898 330186 417134
rect 330422 416898 339186 417134
rect 339422 416898 348186 417134
rect 348422 416898 350748 417134
rect 350984 416898 352400 417134
rect 352636 416898 353206 417134
rect 353442 416898 362206 417134
rect 362442 416898 371206 417134
rect 371442 416898 380206 417134
rect 380442 416898 389206 417134
rect 389442 416898 391768 417134
rect 392004 416898 392420 417134
rect 392656 416898 393226 417134
rect 393462 416898 402226 417134
rect 402462 416898 411226 417134
rect 411462 416898 420226 417134
rect 420462 416898 429226 417134
rect 429462 416898 431788 417134
rect 432024 416898 432440 417134
rect 432676 416898 433246 417134
rect 433482 416898 439792 417134
rect 440028 416898 457010 417134
rect 457246 416898 462842 417134
rect 463078 416898 471028 417134
rect 471264 416898 480028 417134
rect 480264 416898 489028 417134
rect 489264 416898 498028 417134
rect 498264 416898 507028 417134
rect 507264 416898 516028 417134
rect 516264 416898 525028 417134
rect 525264 416898 534028 417134
rect 534264 416898 543028 417134
rect 543264 416898 552028 417134
rect 552264 416898 561028 417134
rect 561264 416898 570028 417134
rect 570264 416898 571450 417134
rect 571686 416898 579470 417134
rect 579706 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 5382 399454
rect 5618 399218 13218 399454
rect 13454 399218 14420 399454
rect 14656 399218 23420 399454
rect 23656 399218 32420 399454
rect 32656 399218 41420 399454
rect 41656 399218 50420 399454
rect 50656 399218 59420 399454
rect 59656 399218 68420 399454
rect 68656 399218 77420 399454
rect 77656 399218 86420 399454
rect 86656 399218 95420 399454
rect 95656 399218 104420 399454
rect 104656 399218 113420 399454
rect 113656 399218 120626 399454
rect 120862 399218 127458 399454
rect 127694 399218 140656 399454
rect 140892 399218 141502 399454
rect 141738 399218 147288 399454
rect 147524 399218 149660 399454
rect 149896 399218 150506 399454
rect 150742 399218 159506 399454
rect 159742 399218 168506 399454
rect 168742 399218 177506 399454
rect 177742 399218 186506 399454
rect 186742 399218 188308 399454
rect 188544 399218 190680 399454
rect 190916 399218 191526 399454
rect 191762 399218 200526 399454
rect 200762 399218 209526 399454
rect 209762 399218 218526 399454
rect 218762 399218 227526 399454
rect 227762 399218 229328 399454
rect 229564 399218 230700 399454
rect 230936 399218 231546 399454
rect 231782 399218 240546 399454
rect 240782 399218 249546 399454
rect 249782 399218 258546 399454
rect 258782 399218 267546 399454
rect 267782 399218 269348 399454
rect 269584 399218 270720 399454
rect 270956 399218 271566 399454
rect 271802 399218 280566 399454
rect 280802 399218 289566 399454
rect 289802 399218 298566 399454
rect 298802 399218 307566 399454
rect 307802 399218 309368 399454
rect 309604 399218 311740 399454
rect 311976 399218 312586 399454
rect 312822 399218 321586 399454
rect 321822 399218 330586 399454
rect 330822 399218 339586 399454
rect 339822 399218 348586 399454
rect 348822 399218 350388 399454
rect 350624 399218 352760 399454
rect 352996 399218 353606 399454
rect 353842 399218 362606 399454
rect 362842 399218 371606 399454
rect 371842 399218 380606 399454
rect 380842 399218 389606 399454
rect 389842 399218 391408 399454
rect 391644 399218 392780 399454
rect 393016 399218 393626 399454
rect 393862 399218 402626 399454
rect 402862 399218 411626 399454
rect 411862 399218 420626 399454
rect 420862 399218 429626 399454
rect 429862 399218 431428 399454
rect 431664 399218 432800 399454
rect 433036 399218 433646 399454
rect 433882 399218 439432 399454
rect 439668 399218 456610 399454
rect 456846 399218 463442 399454
rect 463678 399218 470648 399454
rect 470884 399218 479648 399454
rect 479884 399218 488648 399454
rect 488884 399218 497648 399454
rect 497884 399218 506648 399454
rect 506884 399218 515648 399454
rect 515884 399218 524648 399454
rect 524884 399218 533648 399454
rect 533884 399218 542648 399454
rect 542884 399218 551648 399454
rect 551884 399218 560648 399454
rect 560884 399218 569648 399454
rect 569884 399218 570850 399454
rect 571086 399218 578670 399454
rect 578906 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 5382 399134
rect 5618 398898 13218 399134
rect 13454 398898 14420 399134
rect 14656 398898 23420 399134
rect 23656 398898 32420 399134
rect 32656 398898 41420 399134
rect 41656 398898 50420 399134
rect 50656 398898 59420 399134
rect 59656 398898 68420 399134
rect 68656 398898 77420 399134
rect 77656 398898 86420 399134
rect 86656 398898 95420 399134
rect 95656 398898 104420 399134
rect 104656 398898 113420 399134
rect 113656 398898 120626 399134
rect 120862 398898 127458 399134
rect 127694 398898 140656 399134
rect 140892 398898 141502 399134
rect 141738 398898 147288 399134
rect 147524 398898 149660 399134
rect 149896 398898 150506 399134
rect 150742 398898 159506 399134
rect 159742 398898 168506 399134
rect 168742 398898 177506 399134
rect 177742 398898 186506 399134
rect 186742 398898 188308 399134
rect 188544 398898 190680 399134
rect 190916 398898 191526 399134
rect 191762 398898 200526 399134
rect 200762 398898 209526 399134
rect 209762 398898 218526 399134
rect 218762 398898 227526 399134
rect 227762 398898 229328 399134
rect 229564 398898 230700 399134
rect 230936 398898 231546 399134
rect 231782 398898 240546 399134
rect 240782 398898 249546 399134
rect 249782 398898 258546 399134
rect 258782 398898 267546 399134
rect 267782 398898 269348 399134
rect 269584 398898 270720 399134
rect 270956 398898 271566 399134
rect 271802 398898 280566 399134
rect 280802 398898 289566 399134
rect 289802 398898 298566 399134
rect 298802 398898 307566 399134
rect 307802 398898 309368 399134
rect 309604 398898 311740 399134
rect 311976 398898 312586 399134
rect 312822 398898 321586 399134
rect 321822 398898 330586 399134
rect 330822 398898 339586 399134
rect 339822 398898 348586 399134
rect 348822 398898 350388 399134
rect 350624 398898 352760 399134
rect 352996 398898 353606 399134
rect 353842 398898 362606 399134
rect 362842 398898 371606 399134
rect 371842 398898 380606 399134
rect 380842 398898 389606 399134
rect 389842 398898 391408 399134
rect 391644 398898 392780 399134
rect 393016 398898 393626 399134
rect 393862 398898 402626 399134
rect 402862 398898 411626 399134
rect 411862 398898 420626 399134
rect 420862 398898 429626 399134
rect 429862 398898 431428 399134
rect 431664 398898 432800 399134
rect 433036 398898 433646 399134
rect 433882 398898 439432 399134
rect 439668 398898 456610 399134
rect 456846 398898 463442 399134
rect 463678 398898 470648 399134
rect 470884 398898 479648 399134
rect 479884 398898 488648 399134
rect 488884 398898 497648 399134
rect 497884 398898 506648 399134
rect 506884 398898 515648 399134
rect 515884 398898 524648 399134
rect 524884 398898 533648 399134
rect 533884 398898 542648 399134
rect 542884 398898 551648 399134
rect 551884 398898 560648 399134
rect 560884 398898 569648 399134
rect 569884 398898 570850 399134
rect 571086 398898 578670 399134
rect 578906 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 4582 381454
rect 4818 381218 127058 381454
rect 127294 381218 140296 381454
rect 140532 381218 141102 381454
rect 141338 381218 147648 381454
rect 147884 381218 149300 381454
rect 149536 381218 150106 381454
rect 150342 381218 159106 381454
rect 159342 381218 168106 381454
rect 168342 381218 177106 381454
rect 177342 381218 186106 381454
rect 186342 381218 188668 381454
rect 188904 381218 190320 381454
rect 190556 381218 191126 381454
rect 191362 381218 200126 381454
rect 200362 381218 209126 381454
rect 209362 381218 218126 381454
rect 218362 381218 227126 381454
rect 227362 381218 229688 381454
rect 229924 381218 230340 381454
rect 230576 381218 231146 381454
rect 231382 381218 240146 381454
rect 240382 381218 249146 381454
rect 249382 381218 258146 381454
rect 258382 381218 267146 381454
rect 267382 381218 269708 381454
rect 269944 381218 270360 381454
rect 270596 381218 271166 381454
rect 271402 381218 280166 381454
rect 280402 381218 289166 381454
rect 289402 381218 298166 381454
rect 298402 381218 307166 381454
rect 307402 381218 309728 381454
rect 309964 381218 311380 381454
rect 311616 381218 312186 381454
rect 312422 381218 321186 381454
rect 321422 381218 330186 381454
rect 330422 381218 339186 381454
rect 339422 381218 348186 381454
rect 348422 381218 350748 381454
rect 350984 381218 352400 381454
rect 352636 381218 353206 381454
rect 353442 381218 362206 381454
rect 362442 381218 371206 381454
rect 371442 381218 380206 381454
rect 380442 381218 389206 381454
rect 389442 381218 391768 381454
rect 392004 381218 392420 381454
rect 392656 381218 393226 381454
rect 393462 381218 402226 381454
rect 402462 381218 411226 381454
rect 411462 381218 420226 381454
rect 420462 381218 429226 381454
rect 429462 381218 431788 381454
rect 432024 381218 432440 381454
rect 432676 381218 433246 381454
rect 433482 381218 439792 381454
rect 440028 381218 457010 381454
rect 457246 381218 579470 381454
rect 579706 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 4582 381134
rect 4818 380898 127058 381134
rect 127294 380898 140296 381134
rect 140532 380898 141102 381134
rect 141338 380898 147648 381134
rect 147884 380898 149300 381134
rect 149536 380898 150106 381134
rect 150342 380898 159106 381134
rect 159342 380898 168106 381134
rect 168342 380898 177106 381134
rect 177342 380898 186106 381134
rect 186342 380898 188668 381134
rect 188904 380898 190320 381134
rect 190556 380898 191126 381134
rect 191362 380898 200126 381134
rect 200362 380898 209126 381134
rect 209362 380898 218126 381134
rect 218362 380898 227126 381134
rect 227362 380898 229688 381134
rect 229924 380898 230340 381134
rect 230576 380898 231146 381134
rect 231382 380898 240146 381134
rect 240382 380898 249146 381134
rect 249382 380898 258146 381134
rect 258382 380898 267146 381134
rect 267382 380898 269708 381134
rect 269944 380898 270360 381134
rect 270596 380898 271166 381134
rect 271402 380898 280166 381134
rect 280402 380898 289166 381134
rect 289402 380898 298166 381134
rect 298402 380898 307166 381134
rect 307402 380898 309728 381134
rect 309964 380898 311380 381134
rect 311616 380898 312186 381134
rect 312422 380898 321186 381134
rect 321422 380898 330186 381134
rect 330422 380898 339186 381134
rect 339422 380898 348186 381134
rect 348422 380898 350748 381134
rect 350984 380898 352400 381134
rect 352636 380898 353206 381134
rect 353442 380898 362206 381134
rect 362442 380898 371206 381134
rect 371442 380898 380206 381134
rect 380442 380898 389206 381134
rect 389442 380898 391768 381134
rect 392004 380898 392420 381134
rect 392656 380898 393226 381134
rect 393462 380898 402226 381134
rect 402462 380898 411226 381134
rect 411462 380898 420226 381134
rect 420462 380898 429226 381134
rect 429462 380898 431788 381134
rect 432024 380898 432440 381134
rect 432676 380898 433246 381134
rect 433482 380898 439792 381134
rect 440028 380898 457010 381134
rect 457246 380898 579470 381134
rect 579706 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 5382 363454
rect 5618 363218 127458 363454
rect 127694 363218 140656 363454
rect 140892 363218 141502 363454
rect 141738 363218 147288 363454
rect 147524 363218 149660 363454
rect 149896 363218 150506 363454
rect 150742 363218 159506 363454
rect 159742 363218 168506 363454
rect 168742 363218 177506 363454
rect 177742 363218 186506 363454
rect 186742 363218 188308 363454
rect 188544 363218 190680 363454
rect 190916 363218 191526 363454
rect 191762 363218 200526 363454
rect 200762 363218 209526 363454
rect 209762 363218 218526 363454
rect 218762 363218 227526 363454
rect 227762 363218 229328 363454
rect 229564 363218 230700 363454
rect 230936 363218 231546 363454
rect 231782 363218 240546 363454
rect 240782 363218 249546 363454
rect 249782 363218 258546 363454
rect 258782 363218 267546 363454
rect 267782 363218 269348 363454
rect 269584 363218 270720 363454
rect 270956 363218 271566 363454
rect 271802 363218 280566 363454
rect 280802 363218 289566 363454
rect 289802 363218 298566 363454
rect 298802 363218 307566 363454
rect 307802 363218 309368 363454
rect 309604 363218 311740 363454
rect 311976 363218 312586 363454
rect 312822 363218 321586 363454
rect 321822 363218 330586 363454
rect 330822 363218 339586 363454
rect 339822 363218 348586 363454
rect 348822 363218 350388 363454
rect 350624 363218 352760 363454
rect 352996 363218 353606 363454
rect 353842 363218 362606 363454
rect 362842 363218 371606 363454
rect 371842 363218 380606 363454
rect 380842 363218 389606 363454
rect 389842 363218 391408 363454
rect 391644 363218 392780 363454
rect 393016 363218 393626 363454
rect 393862 363218 402626 363454
rect 402862 363218 411626 363454
rect 411862 363218 420626 363454
rect 420862 363218 429626 363454
rect 429862 363218 431428 363454
rect 431664 363218 432800 363454
rect 433036 363218 433646 363454
rect 433882 363218 439432 363454
rect 439668 363218 456610 363454
rect 456846 363218 578670 363454
rect 578906 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 5382 363134
rect 5618 362898 127458 363134
rect 127694 362898 140656 363134
rect 140892 362898 141502 363134
rect 141738 362898 147288 363134
rect 147524 362898 149660 363134
rect 149896 362898 150506 363134
rect 150742 362898 159506 363134
rect 159742 362898 168506 363134
rect 168742 362898 177506 363134
rect 177742 362898 186506 363134
rect 186742 362898 188308 363134
rect 188544 362898 190680 363134
rect 190916 362898 191526 363134
rect 191762 362898 200526 363134
rect 200762 362898 209526 363134
rect 209762 362898 218526 363134
rect 218762 362898 227526 363134
rect 227762 362898 229328 363134
rect 229564 362898 230700 363134
rect 230936 362898 231546 363134
rect 231782 362898 240546 363134
rect 240782 362898 249546 363134
rect 249782 362898 258546 363134
rect 258782 362898 267546 363134
rect 267782 362898 269348 363134
rect 269584 362898 270720 363134
rect 270956 362898 271566 363134
rect 271802 362898 280566 363134
rect 280802 362898 289566 363134
rect 289802 362898 298566 363134
rect 298802 362898 307566 363134
rect 307802 362898 309368 363134
rect 309604 362898 311740 363134
rect 311976 362898 312586 363134
rect 312822 362898 321586 363134
rect 321822 362898 330586 363134
rect 330822 362898 339586 363134
rect 339822 362898 348586 363134
rect 348822 362898 350388 363134
rect 350624 362898 352760 363134
rect 352996 362898 353606 363134
rect 353842 362898 362606 363134
rect 362842 362898 371606 363134
rect 371842 362898 380606 363134
rect 380842 362898 389606 363134
rect 389842 362898 391408 363134
rect 391644 362898 392780 363134
rect 393016 362898 393626 363134
rect 393862 362898 402626 363134
rect 402862 362898 411626 363134
rect 411862 362898 420626 363134
rect 420862 362898 429626 363134
rect 429862 362898 431428 363134
rect 431664 362898 432800 363134
rect 433036 362898 433646 363134
rect 433882 362898 439432 363134
rect 439668 362898 456610 363134
rect 456846 362898 578670 363134
rect 578906 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 4582 345454
rect 4818 345218 127058 345454
rect 127294 345218 140296 345454
rect 140532 345218 141102 345454
rect 141338 345218 147648 345454
rect 147884 345218 149300 345454
rect 149536 345218 150106 345454
rect 150342 345218 159106 345454
rect 159342 345218 168106 345454
rect 168342 345218 177106 345454
rect 177342 345218 186106 345454
rect 186342 345218 188668 345454
rect 188904 345218 190320 345454
rect 190556 345218 191126 345454
rect 191362 345218 200126 345454
rect 200362 345218 209126 345454
rect 209362 345218 218126 345454
rect 218362 345218 227126 345454
rect 227362 345218 229688 345454
rect 229924 345218 230340 345454
rect 230576 345218 231146 345454
rect 231382 345218 240146 345454
rect 240382 345218 249146 345454
rect 249382 345218 258146 345454
rect 258382 345218 267146 345454
rect 267382 345218 269708 345454
rect 269944 345218 270360 345454
rect 270596 345218 271166 345454
rect 271402 345218 280166 345454
rect 280402 345218 289166 345454
rect 289402 345218 298166 345454
rect 298402 345218 307166 345454
rect 307402 345218 309728 345454
rect 309964 345218 311380 345454
rect 311616 345218 312186 345454
rect 312422 345218 321186 345454
rect 321422 345218 330186 345454
rect 330422 345218 339186 345454
rect 339422 345218 348186 345454
rect 348422 345218 350748 345454
rect 350984 345218 352400 345454
rect 352636 345218 353206 345454
rect 353442 345218 362206 345454
rect 362442 345218 371206 345454
rect 371442 345218 380206 345454
rect 380442 345218 389206 345454
rect 389442 345218 391768 345454
rect 392004 345218 392420 345454
rect 392656 345218 393226 345454
rect 393462 345218 402226 345454
rect 402462 345218 411226 345454
rect 411462 345218 420226 345454
rect 420462 345218 429226 345454
rect 429462 345218 431788 345454
rect 432024 345218 432440 345454
rect 432676 345218 433246 345454
rect 433482 345218 439792 345454
rect 440028 345218 457010 345454
rect 457246 345218 579470 345454
rect 579706 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 4582 345134
rect 4818 344898 127058 345134
rect 127294 344898 140296 345134
rect 140532 344898 141102 345134
rect 141338 344898 147648 345134
rect 147884 344898 149300 345134
rect 149536 344898 150106 345134
rect 150342 344898 159106 345134
rect 159342 344898 168106 345134
rect 168342 344898 177106 345134
rect 177342 344898 186106 345134
rect 186342 344898 188668 345134
rect 188904 344898 190320 345134
rect 190556 344898 191126 345134
rect 191362 344898 200126 345134
rect 200362 344898 209126 345134
rect 209362 344898 218126 345134
rect 218362 344898 227126 345134
rect 227362 344898 229688 345134
rect 229924 344898 230340 345134
rect 230576 344898 231146 345134
rect 231382 344898 240146 345134
rect 240382 344898 249146 345134
rect 249382 344898 258146 345134
rect 258382 344898 267146 345134
rect 267382 344898 269708 345134
rect 269944 344898 270360 345134
rect 270596 344898 271166 345134
rect 271402 344898 280166 345134
rect 280402 344898 289166 345134
rect 289402 344898 298166 345134
rect 298402 344898 307166 345134
rect 307402 344898 309728 345134
rect 309964 344898 311380 345134
rect 311616 344898 312186 345134
rect 312422 344898 321186 345134
rect 321422 344898 330186 345134
rect 330422 344898 339186 345134
rect 339422 344898 348186 345134
rect 348422 344898 350748 345134
rect 350984 344898 352400 345134
rect 352636 344898 353206 345134
rect 353442 344898 362206 345134
rect 362442 344898 371206 345134
rect 371442 344898 380206 345134
rect 380442 344898 389206 345134
rect 389442 344898 391768 345134
rect 392004 344898 392420 345134
rect 392656 344898 393226 345134
rect 393462 344898 402226 345134
rect 402462 344898 411226 345134
rect 411462 344898 420226 345134
rect 420462 344898 429226 345134
rect 429462 344898 431788 345134
rect 432024 344898 432440 345134
rect 432676 344898 433246 345134
rect 433482 344898 439792 345134
rect 440028 344898 457010 345134
rect 457246 344898 579470 345134
rect 579706 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 5382 327454
rect 5618 327218 127458 327454
rect 127694 327218 140656 327454
rect 140892 327218 141502 327454
rect 141738 327218 147288 327454
rect 147524 327218 149660 327454
rect 149896 327218 150506 327454
rect 150742 327218 159506 327454
rect 159742 327218 168506 327454
rect 168742 327218 177506 327454
rect 177742 327218 186506 327454
rect 186742 327218 188308 327454
rect 188544 327218 189768 327454
rect 190004 327218 190680 327454
rect 190916 327218 191526 327454
rect 191762 327218 200526 327454
rect 200762 327218 209526 327454
rect 209762 327218 218526 327454
rect 218762 327218 227526 327454
rect 227762 327218 229328 327454
rect 229564 327218 230700 327454
rect 230936 327218 231546 327454
rect 231782 327218 240546 327454
rect 240782 327218 249546 327454
rect 249782 327218 258546 327454
rect 258782 327218 267546 327454
rect 267782 327218 269348 327454
rect 269584 327218 270720 327454
rect 270956 327218 271566 327454
rect 271802 327218 280566 327454
rect 280802 327218 289566 327454
rect 289802 327218 298566 327454
rect 298802 327218 307566 327454
rect 307802 327218 309368 327454
rect 309604 327218 311740 327454
rect 311976 327218 312586 327454
rect 312822 327218 321586 327454
rect 321822 327218 330586 327454
rect 330822 327218 339586 327454
rect 339822 327218 348586 327454
rect 348822 327218 350388 327454
rect 350624 327218 352760 327454
rect 352996 327218 353606 327454
rect 353842 327218 362606 327454
rect 362842 327218 371606 327454
rect 371842 327218 380606 327454
rect 380842 327218 389606 327454
rect 389842 327218 391408 327454
rect 391644 327218 392780 327454
rect 393016 327218 393626 327454
rect 393862 327218 402626 327454
rect 402862 327218 411626 327454
rect 411862 327218 420626 327454
rect 420862 327218 429626 327454
rect 429862 327218 431428 327454
rect 431664 327218 432800 327454
rect 433036 327218 433646 327454
rect 433882 327218 439432 327454
rect 439668 327218 456610 327454
rect 456846 327218 578670 327454
rect 578906 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 5382 327134
rect 5618 326898 127458 327134
rect 127694 326898 140656 327134
rect 140892 326898 141502 327134
rect 141738 326898 147288 327134
rect 147524 326898 149660 327134
rect 149896 326898 150506 327134
rect 150742 326898 159506 327134
rect 159742 326898 168506 327134
rect 168742 326898 177506 327134
rect 177742 326898 186506 327134
rect 186742 326898 188308 327134
rect 188544 326898 189768 327134
rect 190004 326898 190680 327134
rect 190916 326898 191526 327134
rect 191762 326898 200526 327134
rect 200762 326898 209526 327134
rect 209762 326898 218526 327134
rect 218762 326898 227526 327134
rect 227762 326898 229328 327134
rect 229564 326898 230700 327134
rect 230936 326898 231546 327134
rect 231782 326898 240546 327134
rect 240782 326898 249546 327134
rect 249782 326898 258546 327134
rect 258782 326898 267546 327134
rect 267782 326898 269348 327134
rect 269584 326898 270720 327134
rect 270956 326898 271566 327134
rect 271802 326898 280566 327134
rect 280802 326898 289566 327134
rect 289802 326898 298566 327134
rect 298802 326898 307566 327134
rect 307802 326898 309368 327134
rect 309604 326898 311740 327134
rect 311976 326898 312586 327134
rect 312822 326898 321586 327134
rect 321822 326898 330586 327134
rect 330822 326898 339586 327134
rect 339822 326898 348586 327134
rect 348822 326898 350388 327134
rect 350624 326898 352760 327134
rect 352996 326898 353606 327134
rect 353842 326898 362606 327134
rect 362842 326898 371606 327134
rect 371842 326898 380606 327134
rect 380842 326898 389606 327134
rect 389842 326898 391408 327134
rect 391644 326898 392780 327134
rect 393016 326898 393626 327134
rect 393862 326898 402626 327134
rect 402862 326898 411626 327134
rect 411862 326898 420626 327134
rect 420862 326898 429626 327134
rect 429862 326898 431428 327134
rect 431664 326898 432800 327134
rect 433036 326898 433646 327134
rect 433882 326898 439432 327134
rect 439668 326898 456610 327134
rect 456846 326898 578670 327134
rect 578906 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 4582 309454
rect 4818 309218 127058 309454
rect 127294 309218 140296 309454
rect 140532 309218 141102 309454
rect 141338 309218 147648 309454
rect 147884 309218 149300 309454
rect 149536 309218 150106 309454
rect 150342 309218 159106 309454
rect 159342 309218 168106 309454
rect 168342 309218 177106 309454
rect 177342 309218 186106 309454
rect 186342 309218 188668 309454
rect 188904 309218 190320 309454
rect 190556 309218 191126 309454
rect 191362 309218 200126 309454
rect 200362 309218 209126 309454
rect 209362 309218 218126 309454
rect 218362 309218 227126 309454
rect 227362 309218 229688 309454
rect 229924 309218 230340 309454
rect 230576 309218 231146 309454
rect 231382 309218 240146 309454
rect 240382 309218 249146 309454
rect 249382 309218 258146 309454
rect 258382 309218 267146 309454
rect 267382 309218 269708 309454
rect 269944 309218 270360 309454
rect 270596 309218 271166 309454
rect 271402 309218 280166 309454
rect 280402 309218 289166 309454
rect 289402 309218 298166 309454
rect 298402 309218 307166 309454
rect 307402 309218 309728 309454
rect 309964 309218 311380 309454
rect 311616 309218 312186 309454
rect 312422 309218 321186 309454
rect 321422 309218 330186 309454
rect 330422 309218 339186 309454
rect 339422 309218 348186 309454
rect 348422 309218 350748 309454
rect 350984 309218 352400 309454
rect 352636 309218 353206 309454
rect 353442 309218 362206 309454
rect 362442 309218 371206 309454
rect 371442 309218 380206 309454
rect 380442 309218 389206 309454
rect 389442 309218 391768 309454
rect 392004 309218 392420 309454
rect 392656 309218 393226 309454
rect 393462 309218 402226 309454
rect 402462 309218 411226 309454
rect 411462 309218 420226 309454
rect 420462 309218 429226 309454
rect 429462 309218 431788 309454
rect 432024 309218 432440 309454
rect 432676 309218 433246 309454
rect 433482 309218 439792 309454
rect 440028 309218 457010 309454
rect 457246 309218 579470 309454
rect 579706 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 4582 309134
rect 4818 308898 127058 309134
rect 127294 308898 140296 309134
rect 140532 308898 141102 309134
rect 141338 308898 147648 309134
rect 147884 308898 149300 309134
rect 149536 308898 150106 309134
rect 150342 308898 159106 309134
rect 159342 308898 168106 309134
rect 168342 308898 177106 309134
rect 177342 308898 186106 309134
rect 186342 308898 188668 309134
rect 188904 308898 190320 309134
rect 190556 308898 191126 309134
rect 191362 308898 200126 309134
rect 200362 308898 209126 309134
rect 209362 308898 218126 309134
rect 218362 308898 227126 309134
rect 227362 308898 229688 309134
rect 229924 308898 230340 309134
rect 230576 308898 231146 309134
rect 231382 308898 240146 309134
rect 240382 308898 249146 309134
rect 249382 308898 258146 309134
rect 258382 308898 267146 309134
rect 267382 308898 269708 309134
rect 269944 308898 270360 309134
rect 270596 308898 271166 309134
rect 271402 308898 280166 309134
rect 280402 308898 289166 309134
rect 289402 308898 298166 309134
rect 298402 308898 307166 309134
rect 307402 308898 309728 309134
rect 309964 308898 311380 309134
rect 311616 308898 312186 309134
rect 312422 308898 321186 309134
rect 321422 308898 330186 309134
rect 330422 308898 339186 309134
rect 339422 308898 348186 309134
rect 348422 308898 350748 309134
rect 350984 308898 352400 309134
rect 352636 308898 353206 309134
rect 353442 308898 362206 309134
rect 362442 308898 371206 309134
rect 371442 308898 380206 309134
rect 380442 308898 389206 309134
rect 389442 308898 391768 309134
rect 392004 308898 392420 309134
rect 392656 308898 393226 309134
rect 393462 308898 402226 309134
rect 402462 308898 411226 309134
rect 411462 308898 420226 309134
rect 420462 308898 429226 309134
rect 429462 308898 431788 309134
rect 432024 308898 432440 309134
rect 432676 308898 433246 309134
rect 433482 308898 439792 309134
rect 440028 308898 457010 309134
rect 457246 308898 579470 309134
rect 579706 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 5382 291454
rect 5618 291218 108640 291454
rect 108876 291218 109486 291454
rect 109722 291218 118486 291454
rect 118722 291218 127486 291454
rect 127722 291218 136486 291454
rect 136722 291218 145486 291454
rect 145722 291218 147288 291454
rect 147524 291218 149660 291454
rect 149896 291218 150506 291454
rect 150742 291218 159506 291454
rect 159742 291218 168506 291454
rect 168742 291218 177506 291454
rect 177742 291218 186506 291454
rect 186742 291218 188308 291454
rect 188544 291218 190680 291454
rect 190916 291218 191526 291454
rect 191762 291218 200526 291454
rect 200762 291218 209526 291454
rect 209762 291218 218526 291454
rect 218762 291218 227526 291454
rect 227762 291218 229328 291454
rect 229564 291218 230700 291454
rect 230936 291218 231546 291454
rect 231782 291218 240546 291454
rect 240782 291218 249546 291454
rect 249782 291218 258546 291454
rect 258782 291218 267546 291454
rect 267782 291218 269348 291454
rect 269584 291218 270720 291454
rect 270956 291218 271566 291454
rect 271802 291218 280566 291454
rect 280802 291218 289566 291454
rect 289802 291218 298566 291454
rect 298802 291218 307566 291454
rect 307802 291218 309368 291454
rect 309604 291218 311740 291454
rect 311976 291218 312586 291454
rect 312822 291218 321586 291454
rect 321822 291218 330586 291454
rect 330822 291218 339586 291454
rect 339822 291218 348586 291454
rect 348822 291218 350388 291454
rect 350624 291218 352760 291454
rect 352996 291218 353606 291454
rect 353842 291218 362606 291454
rect 362842 291218 371606 291454
rect 371842 291218 380606 291454
rect 380842 291218 389606 291454
rect 389842 291218 391408 291454
rect 391644 291218 392780 291454
rect 393016 291218 393626 291454
rect 393862 291218 402626 291454
rect 402862 291218 411626 291454
rect 411862 291218 420626 291454
rect 420862 291218 429626 291454
rect 429862 291218 431428 291454
rect 431664 291218 432800 291454
rect 433036 291218 433646 291454
rect 433882 291218 442646 291454
rect 442882 291218 451646 291454
rect 451882 291218 460646 291454
rect 460882 291218 469646 291454
rect 469882 291218 471448 291454
rect 471684 291218 578670 291454
rect 578906 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 5382 291134
rect 5618 290898 108640 291134
rect 108876 290898 109486 291134
rect 109722 290898 118486 291134
rect 118722 290898 127486 291134
rect 127722 290898 136486 291134
rect 136722 290898 145486 291134
rect 145722 290898 147288 291134
rect 147524 290898 149660 291134
rect 149896 290898 150506 291134
rect 150742 290898 159506 291134
rect 159742 290898 168506 291134
rect 168742 290898 177506 291134
rect 177742 290898 186506 291134
rect 186742 290898 188308 291134
rect 188544 290898 190680 291134
rect 190916 290898 191526 291134
rect 191762 290898 200526 291134
rect 200762 290898 209526 291134
rect 209762 290898 218526 291134
rect 218762 290898 227526 291134
rect 227762 290898 229328 291134
rect 229564 290898 230700 291134
rect 230936 290898 231546 291134
rect 231782 290898 240546 291134
rect 240782 290898 249546 291134
rect 249782 290898 258546 291134
rect 258782 290898 267546 291134
rect 267782 290898 269348 291134
rect 269584 290898 270720 291134
rect 270956 290898 271566 291134
rect 271802 290898 280566 291134
rect 280802 290898 289566 291134
rect 289802 290898 298566 291134
rect 298802 290898 307566 291134
rect 307802 290898 309368 291134
rect 309604 290898 311740 291134
rect 311976 290898 312586 291134
rect 312822 290898 321586 291134
rect 321822 290898 330586 291134
rect 330822 290898 339586 291134
rect 339822 290898 348586 291134
rect 348822 290898 350388 291134
rect 350624 290898 352760 291134
rect 352996 290898 353606 291134
rect 353842 290898 362606 291134
rect 362842 290898 371606 291134
rect 371842 290898 380606 291134
rect 380842 290898 389606 291134
rect 389842 290898 391408 291134
rect 391644 290898 392780 291134
rect 393016 290898 393626 291134
rect 393862 290898 402626 291134
rect 402862 290898 411626 291134
rect 411862 290898 420626 291134
rect 420862 290898 429626 291134
rect 429862 290898 431428 291134
rect 431664 290898 432800 291134
rect 433036 290898 433646 291134
rect 433882 290898 442646 291134
rect 442882 290898 451646 291134
rect 451882 290898 460646 291134
rect 460882 290898 469646 291134
rect 469882 290898 471448 291134
rect 471684 290898 578670 291134
rect 578906 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 4582 273454
rect 4818 273218 108280 273454
rect 108516 273218 109086 273454
rect 109322 273218 118086 273454
rect 118322 273218 127086 273454
rect 127322 273218 136086 273454
rect 136322 273218 145086 273454
rect 145322 273218 147648 273454
rect 147884 273218 148782 273454
rect 149018 273218 149300 273454
rect 149536 273218 150106 273454
rect 150342 273218 159106 273454
rect 159342 273218 168106 273454
rect 168342 273218 177106 273454
rect 177342 273218 186106 273454
rect 186342 273218 188668 273454
rect 188904 273218 189216 273454
rect 189452 273218 190320 273454
rect 190556 273218 191126 273454
rect 191362 273218 200126 273454
rect 200362 273218 209126 273454
rect 209362 273218 218126 273454
rect 218362 273218 227126 273454
rect 227362 273218 229688 273454
rect 229924 273218 230340 273454
rect 230576 273218 231146 273454
rect 231382 273218 240146 273454
rect 240382 273218 249146 273454
rect 249382 273218 258146 273454
rect 258382 273218 267146 273454
rect 267382 273218 269708 273454
rect 269944 273218 270360 273454
rect 270596 273218 271166 273454
rect 271402 273218 280166 273454
rect 280402 273218 289166 273454
rect 289402 273218 298166 273454
rect 298402 273218 307166 273454
rect 307402 273218 309728 273454
rect 309964 273218 310840 273454
rect 311076 273218 311380 273454
rect 311616 273218 312186 273454
rect 312422 273218 321186 273454
rect 321422 273218 330186 273454
rect 330422 273218 339186 273454
rect 339422 273218 348186 273454
rect 348422 273218 350748 273454
rect 350984 273218 351320 273454
rect 351556 273218 352400 273454
rect 352636 273218 353206 273454
rect 353442 273218 362206 273454
rect 362442 273218 371206 273454
rect 371442 273218 380206 273454
rect 380442 273218 389206 273454
rect 389442 273218 391768 273454
rect 392004 273218 392420 273454
rect 392656 273218 393226 273454
rect 393462 273218 402226 273454
rect 402462 273218 411226 273454
rect 411462 273218 420226 273454
rect 420462 273218 429226 273454
rect 429462 273218 431788 273454
rect 432024 273218 432440 273454
rect 432676 273218 433246 273454
rect 433482 273218 442246 273454
rect 442482 273218 451246 273454
rect 451482 273218 460246 273454
rect 460482 273218 469246 273454
rect 469482 273218 471808 273454
rect 472044 273218 579470 273454
rect 579706 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 4582 273134
rect 4818 272898 108280 273134
rect 108516 272898 109086 273134
rect 109322 272898 118086 273134
rect 118322 272898 127086 273134
rect 127322 272898 136086 273134
rect 136322 272898 145086 273134
rect 145322 272898 147648 273134
rect 147884 272898 148782 273134
rect 149018 272898 149300 273134
rect 149536 272898 150106 273134
rect 150342 272898 159106 273134
rect 159342 272898 168106 273134
rect 168342 272898 177106 273134
rect 177342 272898 186106 273134
rect 186342 272898 188668 273134
rect 188904 272898 189216 273134
rect 189452 272898 190320 273134
rect 190556 272898 191126 273134
rect 191362 272898 200126 273134
rect 200362 272898 209126 273134
rect 209362 272898 218126 273134
rect 218362 272898 227126 273134
rect 227362 272898 229688 273134
rect 229924 272898 230340 273134
rect 230576 272898 231146 273134
rect 231382 272898 240146 273134
rect 240382 272898 249146 273134
rect 249382 272898 258146 273134
rect 258382 272898 267146 273134
rect 267382 272898 269708 273134
rect 269944 272898 270360 273134
rect 270596 272898 271166 273134
rect 271402 272898 280166 273134
rect 280402 272898 289166 273134
rect 289402 272898 298166 273134
rect 298402 272898 307166 273134
rect 307402 272898 309728 273134
rect 309964 272898 310840 273134
rect 311076 272898 311380 273134
rect 311616 272898 312186 273134
rect 312422 272898 321186 273134
rect 321422 272898 330186 273134
rect 330422 272898 339186 273134
rect 339422 272898 348186 273134
rect 348422 272898 350748 273134
rect 350984 272898 351320 273134
rect 351556 272898 352400 273134
rect 352636 272898 353206 273134
rect 353442 272898 362206 273134
rect 362442 272898 371206 273134
rect 371442 272898 380206 273134
rect 380442 272898 389206 273134
rect 389442 272898 391768 273134
rect 392004 272898 392420 273134
rect 392656 272898 393226 273134
rect 393462 272898 402226 273134
rect 402462 272898 411226 273134
rect 411462 272898 420226 273134
rect 420462 272898 429226 273134
rect 429462 272898 431788 273134
rect 432024 272898 432440 273134
rect 432676 272898 433246 273134
rect 433482 272898 442246 273134
rect 442482 272898 451246 273134
rect 451482 272898 460246 273134
rect 460482 272898 469246 273134
rect 469482 272898 471808 273134
rect 472044 272898 579470 273134
rect 579706 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 5382 255454
rect 5618 255218 12592 255454
rect 12828 255218 13438 255454
rect 13674 255218 22438 255454
rect 22674 255218 27228 255454
rect 27464 255218 28600 255454
rect 28836 255218 29446 255454
rect 29682 255218 38446 255454
rect 38682 255218 47446 255454
rect 47682 255218 56446 255454
rect 56682 255218 65446 255454
rect 65682 255218 67248 255454
rect 67484 255218 68620 255454
rect 68856 255218 69466 255454
rect 69702 255218 78466 255454
rect 78702 255218 87466 255454
rect 87702 255218 96466 255454
rect 96702 255218 105466 255454
rect 105702 255218 107268 255454
rect 107504 255218 108640 255454
rect 108876 255218 109486 255454
rect 109722 255218 118486 255454
rect 118722 255218 127486 255454
rect 127722 255218 136486 255454
rect 136722 255218 145486 255454
rect 145722 255218 147288 255454
rect 147524 255218 149660 255454
rect 149896 255218 150506 255454
rect 150742 255218 159506 255454
rect 159742 255218 168506 255454
rect 168742 255218 177506 255454
rect 177742 255218 186506 255454
rect 186742 255218 188308 255454
rect 188544 255218 190680 255454
rect 190916 255218 191526 255454
rect 191762 255218 200526 255454
rect 200762 255218 209526 255454
rect 209762 255218 218526 255454
rect 218762 255218 227526 255454
rect 227762 255218 229328 255454
rect 229564 255218 230700 255454
rect 230936 255218 231546 255454
rect 231782 255218 240546 255454
rect 240782 255218 249546 255454
rect 249782 255218 258546 255454
rect 258782 255218 267546 255454
rect 267782 255218 269348 255454
rect 269584 255218 270720 255454
rect 270956 255218 271566 255454
rect 271802 255218 280566 255454
rect 280802 255218 289566 255454
rect 289802 255218 298566 255454
rect 298802 255218 307566 255454
rect 307802 255218 309368 255454
rect 309604 255218 311740 255454
rect 311976 255218 312586 255454
rect 312822 255218 321586 255454
rect 321822 255218 330586 255454
rect 330822 255218 339586 255454
rect 339822 255218 348586 255454
rect 348822 255218 350388 255454
rect 350624 255218 352760 255454
rect 352996 255218 353606 255454
rect 353842 255218 362606 255454
rect 362842 255218 371606 255454
rect 371842 255218 380606 255454
rect 380842 255218 389606 255454
rect 389842 255218 391408 255454
rect 391644 255218 392780 255454
rect 393016 255218 393626 255454
rect 393862 255218 402626 255454
rect 402862 255218 411626 255454
rect 411862 255218 420626 255454
rect 420862 255218 429626 255454
rect 429862 255218 431428 255454
rect 431664 255218 432800 255454
rect 433036 255218 433646 255454
rect 433882 255218 442646 255454
rect 442882 255218 451646 255454
rect 451882 255218 460646 255454
rect 460882 255218 469646 255454
rect 469882 255218 471448 255454
rect 471684 255218 472820 255454
rect 473056 255218 473666 255454
rect 473902 255218 482666 255454
rect 482902 255218 491666 255454
rect 491902 255218 500666 255454
rect 500902 255218 509666 255454
rect 509902 255218 511468 255454
rect 511704 255218 512840 255454
rect 513076 255218 513686 255454
rect 513922 255218 522686 255454
rect 522922 255218 531686 255454
rect 531922 255218 540686 255454
rect 540922 255218 549686 255454
rect 549922 255218 551488 255454
rect 551724 255218 552860 255454
rect 553096 255218 553706 255454
rect 553942 255218 562706 255454
rect 562942 255218 571706 255454
rect 571942 255218 573476 255454
rect 573712 255218 578670 255454
rect 578906 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 5382 255134
rect 5618 254898 12592 255134
rect 12828 254898 13438 255134
rect 13674 254898 22438 255134
rect 22674 254898 27228 255134
rect 27464 254898 28600 255134
rect 28836 254898 29446 255134
rect 29682 254898 38446 255134
rect 38682 254898 47446 255134
rect 47682 254898 56446 255134
rect 56682 254898 65446 255134
rect 65682 254898 67248 255134
rect 67484 254898 68620 255134
rect 68856 254898 69466 255134
rect 69702 254898 78466 255134
rect 78702 254898 87466 255134
rect 87702 254898 96466 255134
rect 96702 254898 105466 255134
rect 105702 254898 107268 255134
rect 107504 254898 108640 255134
rect 108876 254898 109486 255134
rect 109722 254898 118486 255134
rect 118722 254898 127486 255134
rect 127722 254898 136486 255134
rect 136722 254898 145486 255134
rect 145722 254898 147288 255134
rect 147524 254898 149660 255134
rect 149896 254898 150506 255134
rect 150742 254898 159506 255134
rect 159742 254898 168506 255134
rect 168742 254898 177506 255134
rect 177742 254898 186506 255134
rect 186742 254898 188308 255134
rect 188544 254898 190680 255134
rect 190916 254898 191526 255134
rect 191762 254898 200526 255134
rect 200762 254898 209526 255134
rect 209762 254898 218526 255134
rect 218762 254898 227526 255134
rect 227762 254898 229328 255134
rect 229564 254898 230700 255134
rect 230936 254898 231546 255134
rect 231782 254898 240546 255134
rect 240782 254898 249546 255134
rect 249782 254898 258546 255134
rect 258782 254898 267546 255134
rect 267782 254898 269348 255134
rect 269584 254898 270720 255134
rect 270956 254898 271566 255134
rect 271802 254898 280566 255134
rect 280802 254898 289566 255134
rect 289802 254898 298566 255134
rect 298802 254898 307566 255134
rect 307802 254898 309368 255134
rect 309604 254898 311740 255134
rect 311976 254898 312586 255134
rect 312822 254898 321586 255134
rect 321822 254898 330586 255134
rect 330822 254898 339586 255134
rect 339822 254898 348586 255134
rect 348822 254898 350388 255134
rect 350624 254898 352760 255134
rect 352996 254898 353606 255134
rect 353842 254898 362606 255134
rect 362842 254898 371606 255134
rect 371842 254898 380606 255134
rect 380842 254898 389606 255134
rect 389842 254898 391408 255134
rect 391644 254898 392780 255134
rect 393016 254898 393626 255134
rect 393862 254898 402626 255134
rect 402862 254898 411626 255134
rect 411862 254898 420626 255134
rect 420862 254898 429626 255134
rect 429862 254898 431428 255134
rect 431664 254898 432800 255134
rect 433036 254898 433646 255134
rect 433882 254898 442646 255134
rect 442882 254898 451646 255134
rect 451882 254898 460646 255134
rect 460882 254898 469646 255134
rect 469882 254898 471448 255134
rect 471684 254898 472820 255134
rect 473056 254898 473666 255134
rect 473902 254898 482666 255134
rect 482902 254898 491666 255134
rect 491902 254898 500666 255134
rect 500902 254898 509666 255134
rect 509902 254898 511468 255134
rect 511704 254898 512840 255134
rect 513076 254898 513686 255134
rect 513922 254898 522686 255134
rect 522922 254898 531686 255134
rect 531922 254898 540686 255134
rect 540922 254898 549686 255134
rect 549922 254898 551488 255134
rect 551724 254898 552860 255134
rect 553096 254898 553706 255134
rect 553942 254898 562706 255134
rect 562942 254898 571706 255134
rect 571942 254898 573476 255134
rect 573712 254898 578670 255134
rect 578906 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 4582 237454
rect 4818 237218 12232 237454
rect 12468 237218 13038 237454
rect 13274 237218 22038 237454
rect 22274 237218 27588 237454
rect 27824 237218 28240 237454
rect 28476 237218 29046 237454
rect 29282 237218 38046 237454
rect 38282 237218 47046 237454
rect 47282 237218 56046 237454
rect 56282 237218 65046 237454
rect 65282 237218 67608 237454
rect 67844 237218 68260 237454
rect 68496 237218 69066 237454
rect 69302 237218 78066 237454
rect 78302 237218 87066 237454
rect 87302 237218 96066 237454
rect 96302 237218 105066 237454
rect 105302 237218 107628 237454
rect 107864 237218 108280 237454
rect 108516 237218 109086 237454
rect 109322 237218 118086 237454
rect 118322 237218 127086 237454
rect 127322 237218 136086 237454
rect 136322 237218 145086 237454
rect 145322 237218 147648 237454
rect 147884 237218 148782 237454
rect 149018 237218 149300 237454
rect 149536 237218 150106 237454
rect 150342 237218 159106 237454
rect 159342 237218 168106 237454
rect 168342 237218 177106 237454
rect 177342 237218 186106 237454
rect 186342 237218 188668 237454
rect 188904 237218 189216 237454
rect 189452 237218 190320 237454
rect 190556 237218 191126 237454
rect 191362 237218 200126 237454
rect 200362 237218 209126 237454
rect 209362 237218 218126 237454
rect 218362 237218 227126 237454
rect 227362 237218 229688 237454
rect 229924 237218 230340 237454
rect 230576 237218 231146 237454
rect 231382 237218 240146 237454
rect 240382 237218 249146 237454
rect 249382 237218 258146 237454
rect 258382 237218 267146 237454
rect 267382 237218 269708 237454
rect 269944 237218 270360 237454
rect 270596 237218 271166 237454
rect 271402 237218 280166 237454
rect 280402 237218 289166 237454
rect 289402 237218 298166 237454
rect 298402 237218 307166 237454
rect 307402 237218 309728 237454
rect 309964 237218 310840 237454
rect 311076 237218 311380 237454
rect 311616 237218 312186 237454
rect 312422 237218 321186 237454
rect 321422 237218 330186 237454
rect 330422 237218 339186 237454
rect 339422 237218 348186 237454
rect 348422 237218 350748 237454
rect 350984 237218 351320 237454
rect 351556 237218 352400 237454
rect 352636 237218 353206 237454
rect 353442 237218 362206 237454
rect 362442 237218 371206 237454
rect 371442 237218 380206 237454
rect 380442 237218 389206 237454
rect 389442 237218 391768 237454
rect 392004 237218 392420 237454
rect 392656 237218 393226 237454
rect 393462 237218 402226 237454
rect 402462 237218 411226 237454
rect 411462 237218 420226 237454
rect 420462 237218 429226 237454
rect 429462 237218 431788 237454
rect 432024 237218 432440 237454
rect 432676 237218 433246 237454
rect 433482 237218 442246 237454
rect 442482 237218 451246 237454
rect 451482 237218 460246 237454
rect 460482 237218 469246 237454
rect 469482 237218 471808 237454
rect 472044 237218 472460 237454
rect 472696 237218 473266 237454
rect 473502 237218 482266 237454
rect 482502 237218 491266 237454
rect 491502 237218 500266 237454
rect 500502 237218 509266 237454
rect 509502 237218 511828 237454
rect 512064 237218 512480 237454
rect 512716 237218 513286 237454
rect 513522 237218 522286 237454
rect 522522 237218 531286 237454
rect 531522 237218 540286 237454
rect 540522 237218 549286 237454
rect 549522 237218 551848 237454
rect 552084 237218 552500 237454
rect 552736 237218 553306 237454
rect 553542 237218 562306 237454
rect 562542 237218 571306 237454
rect 571542 237218 573836 237454
rect 574072 237218 579470 237454
rect 579706 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 4582 237134
rect 4818 236898 12232 237134
rect 12468 236898 13038 237134
rect 13274 236898 22038 237134
rect 22274 236898 27588 237134
rect 27824 236898 28240 237134
rect 28476 236898 29046 237134
rect 29282 236898 38046 237134
rect 38282 236898 47046 237134
rect 47282 236898 56046 237134
rect 56282 236898 65046 237134
rect 65282 236898 67608 237134
rect 67844 236898 68260 237134
rect 68496 236898 69066 237134
rect 69302 236898 78066 237134
rect 78302 236898 87066 237134
rect 87302 236898 96066 237134
rect 96302 236898 105066 237134
rect 105302 236898 107628 237134
rect 107864 236898 108280 237134
rect 108516 236898 109086 237134
rect 109322 236898 118086 237134
rect 118322 236898 127086 237134
rect 127322 236898 136086 237134
rect 136322 236898 145086 237134
rect 145322 236898 147648 237134
rect 147884 236898 148782 237134
rect 149018 236898 149300 237134
rect 149536 236898 150106 237134
rect 150342 236898 159106 237134
rect 159342 236898 168106 237134
rect 168342 236898 177106 237134
rect 177342 236898 186106 237134
rect 186342 236898 188668 237134
rect 188904 236898 189216 237134
rect 189452 236898 190320 237134
rect 190556 236898 191126 237134
rect 191362 236898 200126 237134
rect 200362 236898 209126 237134
rect 209362 236898 218126 237134
rect 218362 236898 227126 237134
rect 227362 236898 229688 237134
rect 229924 236898 230340 237134
rect 230576 236898 231146 237134
rect 231382 236898 240146 237134
rect 240382 236898 249146 237134
rect 249382 236898 258146 237134
rect 258382 236898 267146 237134
rect 267382 236898 269708 237134
rect 269944 236898 270360 237134
rect 270596 236898 271166 237134
rect 271402 236898 280166 237134
rect 280402 236898 289166 237134
rect 289402 236898 298166 237134
rect 298402 236898 307166 237134
rect 307402 236898 309728 237134
rect 309964 236898 310840 237134
rect 311076 236898 311380 237134
rect 311616 236898 312186 237134
rect 312422 236898 321186 237134
rect 321422 236898 330186 237134
rect 330422 236898 339186 237134
rect 339422 236898 348186 237134
rect 348422 236898 350748 237134
rect 350984 236898 351320 237134
rect 351556 236898 352400 237134
rect 352636 236898 353206 237134
rect 353442 236898 362206 237134
rect 362442 236898 371206 237134
rect 371442 236898 380206 237134
rect 380442 236898 389206 237134
rect 389442 236898 391768 237134
rect 392004 236898 392420 237134
rect 392656 236898 393226 237134
rect 393462 236898 402226 237134
rect 402462 236898 411226 237134
rect 411462 236898 420226 237134
rect 420462 236898 429226 237134
rect 429462 236898 431788 237134
rect 432024 236898 432440 237134
rect 432676 236898 433246 237134
rect 433482 236898 442246 237134
rect 442482 236898 451246 237134
rect 451482 236898 460246 237134
rect 460482 236898 469246 237134
rect 469482 236898 471808 237134
rect 472044 236898 472460 237134
rect 472696 236898 473266 237134
rect 473502 236898 482266 237134
rect 482502 236898 491266 237134
rect 491502 236898 500266 237134
rect 500502 236898 509266 237134
rect 509502 236898 511828 237134
rect 512064 236898 512480 237134
rect 512716 236898 513286 237134
rect 513522 236898 522286 237134
rect 522522 236898 531286 237134
rect 531522 236898 540286 237134
rect 540522 236898 549286 237134
rect 549522 236898 551848 237134
rect 552084 236898 552500 237134
rect 552736 236898 553306 237134
rect 553542 236898 562306 237134
rect 562542 236898 571306 237134
rect 571542 236898 573836 237134
rect 574072 236898 579470 237134
rect 579706 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 5382 219454
rect 5618 219218 12592 219454
rect 12828 219218 13438 219454
rect 13674 219218 22438 219454
rect 22674 219218 27228 219454
rect 27464 219218 28600 219454
rect 28836 219218 29446 219454
rect 29682 219218 38446 219454
rect 38682 219218 47446 219454
rect 47682 219218 56446 219454
rect 56682 219218 65446 219454
rect 65682 219218 67248 219454
rect 67484 219218 68620 219454
rect 68856 219218 69466 219454
rect 69702 219218 78466 219454
rect 78702 219218 87466 219454
rect 87702 219218 96466 219454
rect 96702 219218 105466 219454
rect 105702 219218 107268 219454
rect 107504 219218 108640 219454
rect 108876 219218 109486 219454
rect 109722 219218 118486 219454
rect 118722 219218 127486 219454
rect 127722 219218 136486 219454
rect 136722 219218 145486 219454
rect 145722 219218 147288 219454
rect 147524 219218 149660 219454
rect 149896 219218 150506 219454
rect 150742 219218 159506 219454
rect 159742 219218 168506 219454
rect 168742 219218 177506 219454
rect 177742 219218 186506 219454
rect 186742 219218 188308 219454
rect 188544 219218 190680 219454
rect 190916 219218 191526 219454
rect 191762 219218 200526 219454
rect 200762 219218 209526 219454
rect 209762 219218 218526 219454
rect 218762 219218 227526 219454
rect 227762 219218 229328 219454
rect 229564 219218 230700 219454
rect 230936 219218 231546 219454
rect 231782 219218 240546 219454
rect 240782 219218 249546 219454
rect 249782 219218 258546 219454
rect 258782 219218 267546 219454
rect 267782 219218 269348 219454
rect 269584 219218 270720 219454
rect 270956 219218 271566 219454
rect 271802 219218 280566 219454
rect 280802 219218 289566 219454
rect 289802 219218 298566 219454
rect 298802 219218 307566 219454
rect 307802 219218 309368 219454
rect 309604 219218 311740 219454
rect 311976 219218 312586 219454
rect 312822 219218 321586 219454
rect 321822 219218 330586 219454
rect 330822 219218 339586 219454
rect 339822 219218 348586 219454
rect 348822 219218 350388 219454
rect 350624 219218 352760 219454
rect 352996 219218 353606 219454
rect 353842 219218 362606 219454
rect 362842 219218 371606 219454
rect 371842 219218 380606 219454
rect 380842 219218 389606 219454
rect 389842 219218 391408 219454
rect 391644 219218 392780 219454
rect 393016 219218 393626 219454
rect 393862 219218 402626 219454
rect 402862 219218 411626 219454
rect 411862 219218 420626 219454
rect 420862 219218 429626 219454
rect 429862 219218 431428 219454
rect 431664 219218 432800 219454
rect 433036 219218 433646 219454
rect 433882 219218 442646 219454
rect 442882 219218 451646 219454
rect 451882 219218 460646 219454
rect 460882 219218 469646 219454
rect 469882 219218 471448 219454
rect 471684 219218 472820 219454
rect 473056 219218 473666 219454
rect 473902 219218 482666 219454
rect 482902 219218 491666 219454
rect 491902 219218 500666 219454
rect 500902 219218 509666 219454
rect 509902 219218 511468 219454
rect 511704 219218 512840 219454
rect 513076 219218 513686 219454
rect 513922 219218 522686 219454
rect 522922 219218 531686 219454
rect 531922 219218 540686 219454
rect 540922 219218 549686 219454
rect 549922 219218 551488 219454
rect 551724 219218 552860 219454
rect 553096 219218 553706 219454
rect 553942 219218 562706 219454
rect 562942 219218 571706 219454
rect 571942 219218 573476 219454
rect 573712 219218 578670 219454
rect 578906 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 5382 219134
rect 5618 218898 12592 219134
rect 12828 218898 13438 219134
rect 13674 218898 22438 219134
rect 22674 218898 27228 219134
rect 27464 218898 28600 219134
rect 28836 218898 29446 219134
rect 29682 218898 38446 219134
rect 38682 218898 47446 219134
rect 47682 218898 56446 219134
rect 56682 218898 65446 219134
rect 65682 218898 67248 219134
rect 67484 218898 68620 219134
rect 68856 218898 69466 219134
rect 69702 218898 78466 219134
rect 78702 218898 87466 219134
rect 87702 218898 96466 219134
rect 96702 218898 105466 219134
rect 105702 218898 107268 219134
rect 107504 218898 108640 219134
rect 108876 218898 109486 219134
rect 109722 218898 118486 219134
rect 118722 218898 127486 219134
rect 127722 218898 136486 219134
rect 136722 218898 145486 219134
rect 145722 218898 147288 219134
rect 147524 218898 149660 219134
rect 149896 218898 150506 219134
rect 150742 218898 159506 219134
rect 159742 218898 168506 219134
rect 168742 218898 177506 219134
rect 177742 218898 186506 219134
rect 186742 218898 188308 219134
rect 188544 218898 190680 219134
rect 190916 218898 191526 219134
rect 191762 218898 200526 219134
rect 200762 218898 209526 219134
rect 209762 218898 218526 219134
rect 218762 218898 227526 219134
rect 227762 218898 229328 219134
rect 229564 218898 230700 219134
rect 230936 218898 231546 219134
rect 231782 218898 240546 219134
rect 240782 218898 249546 219134
rect 249782 218898 258546 219134
rect 258782 218898 267546 219134
rect 267782 218898 269348 219134
rect 269584 218898 270720 219134
rect 270956 218898 271566 219134
rect 271802 218898 280566 219134
rect 280802 218898 289566 219134
rect 289802 218898 298566 219134
rect 298802 218898 307566 219134
rect 307802 218898 309368 219134
rect 309604 218898 311740 219134
rect 311976 218898 312586 219134
rect 312822 218898 321586 219134
rect 321822 218898 330586 219134
rect 330822 218898 339586 219134
rect 339822 218898 348586 219134
rect 348822 218898 350388 219134
rect 350624 218898 352760 219134
rect 352996 218898 353606 219134
rect 353842 218898 362606 219134
rect 362842 218898 371606 219134
rect 371842 218898 380606 219134
rect 380842 218898 389606 219134
rect 389842 218898 391408 219134
rect 391644 218898 392780 219134
rect 393016 218898 393626 219134
rect 393862 218898 402626 219134
rect 402862 218898 411626 219134
rect 411862 218898 420626 219134
rect 420862 218898 429626 219134
rect 429862 218898 431428 219134
rect 431664 218898 432800 219134
rect 433036 218898 433646 219134
rect 433882 218898 442646 219134
rect 442882 218898 451646 219134
rect 451882 218898 460646 219134
rect 460882 218898 469646 219134
rect 469882 218898 471448 219134
rect 471684 218898 472820 219134
rect 473056 218898 473666 219134
rect 473902 218898 482666 219134
rect 482902 218898 491666 219134
rect 491902 218898 500666 219134
rect 500902 218898 509666 219134
rect 509902 218898 511468 219134
rect 511704 218898 512840 219134
rect 513076 218898 513686 219134
rect 513922 218898 522686 219134
rect 522922 218898 531686 219134
rect 531922 218898 540686 219134
rect 540922 218898 549686 219134
rect 549922 218898 551488 219134
rect 551724 218898 552860 219134
rect 553096 218898 553706 219134
rect 553942 218898 562706 219134
rect 562942 218898 571706 219134
rect 571942 218898 573476 219134
rect 573712 218898 578670 219134
rect 578906 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 4582 201454
rect 4818 201218 12232 201454
rect 12468 201218 13038 201454
rect 13274 201218 22038 201454
rect 22274 201218 27588 201454
rect 27824 201218 28240 201454
rect 28476 201218 29046 201454
rect 29282 201218 38046 201454
rect 38282 201218 47046 201454
rect 47282 201218 56046 201454
rect 56282 201218 65046 201454
rect 65282 201218 67608 201454
rect 67844 201218 68260 201454
rect 68496 201218 69066 201454
rect 69302 201218 78066 201454
rect 78302 201218 87066 201454
rect 87302 201218 96066 201454
rect 96302 201218 105066 201454
rect 105302 201218 107628 201454
rect 107864 201218 108280 201454
rect 108516 201218 109086 201454
rect 109322 201218 118086 201454
rect 118322 201218 127086 201454
rect 127322 201218 136086 201454
rect 136322 201218 145086 201454
rect 145322 201218 147648 201454
rect 147884 201218 149300 201454
rect 149536 201218 150106 201454
rect 150342 201218 159106 201454
rect 159342 201218 168106 201454
rect 168342 201218 177106 201454
rect 177342 201218 186106 201454
rect 186342 201218 188668 201454
rect 188904 201218 190320 201454
rect 190556 201218 191126 201454
rect 191362 201218 200126 201454
rect 200362 201218 209126 201454
rect 209362 201218 218126 201454
rect 218362 201218 227126 201454
rect 227362 201218 229688 201454
rect 229924 201218 230340 201454
rect 230576 201218 231146 201454
rect 231382 201218 240146 201454
rect 240382 201218 249146 201454
rect 249382 201218 258146 201454
rect 258382 201218 267146 201454
rect 267382 201218 269708 201454
rect 269944 201218 270360 201454
rect 270596 201218 271166 201454
rect 271402 201218 280166 201454
rect 280402 201218 289166 201454
rect 289402 201218 298166 201454
rect 298402 201218 307166 201454
rect 307402 201218 309728 201454
rect 309964 201218 311380 201454
rect 311616 201218 312186 201454
rect 312422 201218 321186 201454
rect 321422 201218 330186 201454
rect 330422 201218 339186 201454
rect 339422 201218 348186 201454
rect 348422 201218 350748 201454
rect 350984 201218 352400 201454
rect 352636 201218 353206 201454
rect 353442 201218 362206 201454
rect 362442 201218 371206 201454
rect 371442 201218 380206 201454
rect 380442 201218 389206 201454
rect 389442 201218 391768 201454
rect 392004 201218 392420 201454
rect 392656 201218 393226 201454
rect 393462 201218 402226 201454
rect 402462 201218 411226 201454
rect 411462 201218 420226 201454
rect 420462 201218 429226 201454
rect 429462 201218 431788 201454
rect 432024 201218 432440 201454
rect 432676 201218 433246 201454
rect 433482 201218 442246 201454
rect 442482 201218 451246 201454
rect 451482 201218 460246 201454
rect 460482 201218 469246 201454
rect 469482 201218 471808 201454
rect 472044 201218 472460 201454
rect 472696 201218 473266 201454
rect 473502 201218 482266 201454
rect 482502 201218 491266 201454
rect 491502 201218 500266 201454
rect 500502 201218 509266 201454
rect 509502 201218 511828 201454
rect 512064 201218 512480 201454
rect 512716 201218 513286 201454
rect 513522 201218 522286 201454
rect 522522 201218 531286 201454
rect 531522 201218 540286 201454
rect 540522 201218 549286 201454
rect 549522 201218 551848 201454
rect 552084 201218 552500 201454
rect 552736 201218 553306 201454
rect 553542 201218 562306 201454
rect 562542 201218 571306 201454
rect 571542 201218 573836 201454
rect 574072 201218 579470 201454
rect 579706 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 4582 201134
rect 4818 200898 12232 201134
rect 12468 200898 13038 201134
rect 13274 200898 22038 201134
rect 22274 200898 27588 201134
rect 27824 200898 28240 201134
rect 28476 200898 29046 201134
rect 29282 200898 38046 201134
rect 38282 200898 47046 201134
rect 47282 200898 56046 201134
rect 56282 200898 65046 201134
rect 65282 200898 67608 201134
rect 67844 200898 68260 201134
rect 68496 200898 69066 201134
rect 69302 200898 78066 201134
rect 78302 200898 87066 201134
rect 87302 200898 96066 201134
rect 96302 200898 105066 201134
rect 105302 200898 107628 201134
rect 107864 200898 108280 201134
rect 108516 200898 109086 201134
rect 109322 200898 118086 201134
rect 118322 200898 127086 201134
rect 127322 200898 136086 201134
rect 136322 200898 145086 201134
rect 145322 200898 147648 201134
rect 147884 200898 149300 201134
rect 149536 200898 150106 201134
rect 150342 200898 159106 201134
rect 159342 200898 168106 201134
rect 168342 200898 177106 201134
rect 177342 200898 186106 201134
rect 186342 200898 188668 201134
rect 188904 200898 190320 201134
rect 190556 200898 191126 201134
rect 191362 200898 200126 201134
rect 200362 200898 209126 201134
rect 209362 200898 218126 201134
rect 218362 200898 227126 201134
rect 227362 200898 229688 201134
rect 229924 200898 230340 201134
rect 230576 200898 231146 201134
rect 231382 200898 240146 201134
rect 240382 200898 249146 201134
rect 249382 200898 258146 201134
rect 258382 200898 267146 201134
rect 267382 200898 269708 201134
rect 269944 200898 270360 201134
rect 270596 200898 271166 201134
rect 271402 200898 280166 201134
rect 280402 200898 289166 201134
rect 289402 200898 298166 201134
rect 298402 200898 307166 201134
rect 307402 200898 309728 201134
rect 309964 200898 311380 201134
rect 311616 200898 312186 201134
rect 312422 200898 321186 201134
rect 321422 200898 330186 201134
rect 330422 200898 339186 201134
rect 339422 200898 348186 201134
rect 348422 200898 350748 201134
rect 350984 200898 352400 201134
rect 352636 200898 353206 201134
rect 353442 200898 362206 201134
rect 362442 200898 371206 201134
rect 371442 200898 380206 201134
rect 380442 200898 389206 201134
rect 389442 200898 391768 201134
rect 392004 200898 392420 201134
rect 392656 200898 393226 201134
rect 393462 200898 402226 201134
rect 402462 200898 411226 201134
rect 411462 200898 420226 201134
rect 420462 200898 429226 201134
rect 429462 200898 431788 201134
rect 432024 200898 432440 201134
rect 432676 200898 433246 201134
rect 433482 200898 442246 201134
rect 442482 200898 451246 201134
rect 451482 200898 460246 201134
rect 460482 200898 469246 201134
rect 469482 200898 471808 201134
rect 472044 200898 472460 201134
rect 472696 200898 473266 201134
rect 473502 200898 482266 201134
rect 482502 200898 491266 201134
rect 491502 200898 500266 201134
rect 500502 200898 509266 201134
rect 509502 200898 511828 201134
rect 512064 200898 512480 201134
rect 512716 200898 513286 201134
rect 513522 200898 522286 201134
rect 522522 200898 531286 201134
rect 531522 200898 540286 201134
rect 540522 200898 549286 201134
rect 549522 200898 551848 201134
rect 552084 200898 552500 201134
rect 552736 200898 553306 201134
rect 553542 200898 562306 201134
rect 562542 200898 571306 201134
rect 571542 200898 573836 201134
rect 574072 200898 579470 201134
rect 579706 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 5382 183454
rect 5618 183218 12592 183454
rect 12828 183218 13438 183454
rect 13674 183218 22438 183454
rect 22674 183218 27228 183454
rect 27464 183218 28600 183454
rect 28836 183218 29446 183454
rect 29682 183218 38446 183454
rect 38682 183218 47446 183454
rect 47682 183218 56446 183454
rect 56682 183218 65446 183454
rect 65682 183218 67248 183454
rect 67484 183218 68620 183454
rect 68856 183218 69466 183454
rect 69702 183218 78466 183454
rect 78702 183218 87466 183454
rect 87702 183218 96466 183454
rect 96702 183218 105466 183454
rect 105702 183218 107268 183454
rect 107504 183218 108640 183454
rect 108876 183218 109486 183454
rect 109722 183218 118486 183454
rect 118722 183218 127486 183454
rect 127722 183218 136486 183454
rect 136722 183218 145486 183454
rect 145722 183218 147288 183454
rect 147524 183218 149660 183454
rect 149896 183218 150506 183454
rect 150742 183218 159506 183454
rect 159742 183218 168506 183454
rect 168742 183218 177506 183454
rect 177742 183218 186506 183454
rect 186742 183218 188308 183454
rect 188544 183218 190680 183454
rect 190916 183218 191526 183454
rect 191762 183218 200526 183454
rect 200762 183218 209526 183454
rect 209762 183218 218526 183454
rect 218762 183218 227526 183454
rect 227762 183218 229328 183454
rect 229564 183218 230700 183454
rect 230936 183218 231546 183454
rect 231782 183218 240546 183454
rect 240782 183218 249546 183454
rect 249782 183218 258546 183454
rect 258782 183218 267546 183454
rect 267782 183218 269348 183454
rect 269584 183218 270720 183454
rect 270956 183218 271566 183454
rect 271802 183218 280566 183454
rect 280802 183218 289566 183454
rect 289802 183218 298566 183454
rect 298802 183218 307566 183454
rect 307802 183218 309368 183454
rect 309604 183218 311740 183454
rect 311976 183218 312586 183454
rect 312822 183218 321586 183454
rect 321822 183218 330586 183454
rect 330822 183218 339586 183454
rect 339822 183218 348586 183454
rect 348822 183218 350388 183454
rect 350624 183218 352760 183454
rect 352996 183218 353606 183454
rect 353842 183218 362606 183454
rect 362842 183218 371606 183454
rect 371842 183218 380606 183454
rect 380842 183218 389606 183454
rect 389842 183218 391408 183454
rect 391644 183218 392780 183454
rect 393016 183218 393626 183454
rect 393862 183218 402626 183454
rect 402862 183218 411626 183454
rect 411862 183218 420626 183454
rect 420862 183218 429626 183454
rect 429862 183218 431428 183454
rect 431664 183218 432800 183454
rect 433036 183218 433646 183454
rect 433882 183218 442646 183454
rect 442882 183218 451646 183454
rect 451882 183218 460646 183454
rect 460882 183218 469646 183454
rect 469882 183218 471448 183454
rect 471684 183218 472820 183454
rect 473056 183218 473666 183454
rect 473902 183218 482666 183454
rect 482902 183218 491666 183454
rect 491902 183218 500666 183454
rect 500902 183218 509666 183454
rect 509902 183218 511468 183454
rect 511704 183218 512840 183454
rect 513076 183218 513686 183454
rect 513922 183218 522686 183454
rect 522922 183218 531686 183454
rect 531922 183218 540686 183454
rect 540922 183218 549686 183454
rect 549922 183218 551488 183454
rect 551724 183218 552860 183454
rect 553096 183218 553706 183454
rect 553942 183218 562706 183454
rect 562942 183218 571706 183454
rect 571942 183218 573476 183454
rect 573712 183218 578670 183454
rect 578906 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 5382 183134
rect 5618 182898 12592 183134
rect 12828 182898 13438 183134
rect 13674 182898 22438 183134
rect 22674 182898 27228 183134
rect 27464 182898 28600 183134
rect 28836 182898 29446 183134
rect 29682 182898 38446 183134
rect 38682 182898 47446 183134
rect 47682 182898 56446 183134
rect 56682 182898 65446 183134
rect 65682 182898 67248 183134
rect 67484 182898 68620 183134
rect 68856 182898 69466 183134
rect 69702 182898 78466 183134
rect 78702 182898 87466 183134
rect 87702 182898 96466 183134
rect 96702 182898 105466 183134
rect 105702 182898 107268 183134
rect 107504 182898 108640 183134
rect 108876 182898 109486 183134
rect 109722 182898 118486 183134
rect 118722 182898 127486 183134
rect 127722 182898 136486 183134
rect 136722 182898 145486 183134
rect 145722 182898 147288 183134
rect 147524 182898 149660 183134
rect 149896 182898 150506 183134
rect 150742 182898 159506 183134
rect 159742 182898 168506 183134
rect 168742 182898 177506 183134
rect 177742 182898 186506 183134
rect 186742 182898 188308 183134
rect 188544 182898 190680 183134
rect 190916 182898 191526 183134
rect 191762 182898 200526 183134
rect 200762 182898 209526 183134
rect 209762 182898 218526 183134
rect 218762 182898 227526 183134
rect 227762 182898 229328 183134
rect 229564 182898 230700 183134
rect 230936 182898 231546 183134
rect 231782 182898 240546 183134
rect 240782 182898 249546 183134
rect 249782 182898 258546 183134
rect 258782 182898 267546 183134
rect 267782 182898 269348 183134
rect 269584 182898 270720 183134
rect 270956 182898 271566 183134
rect 271802 182898 280566 183134
rect 280802 182898 289566 183134
rect 289802 182898 298566 183134
rect 298802 182898 307566 183134
rect 307802 182898 309368 183134
rect 309604 182898 311740 183134
rect 311976 182898 312586 183134
rect 312822 182898 321586 183134
rect 321822 182898 330586 183134
rect 330822 182898 339586 183134
rect 339822 182898 348586 183134
rect 348822 182898 350388 183134
rect 350624 182898 352760 183134
rect 352996 182898 353606 183134
rect 353842 182898 362606 183134
rect 362842 182898 371606 183134
rect 371842 182898 380606 183134
rect 380842 182898 389606 183134
rect 389842 182898 391408 183134
rect 391644 182898 392780 183134
rect 393016 182898 393626 183134
rect 393862 182898 402626 183134
rect 402862 182898 411626 183134
rect 411862 182898 420626 183134
rect 420862 182898 429626 183134
rect 429862 182898 431428 183134
rect 431664 182898 432800 183134
rect 433036 182898 433646 183134
rect 433882 182898 442646 183134
rect 442882 182898 451646 183134
rect 451882 182898 460646 183134
rect 460882 182898 469646 183134
rect 469882 182898 471448 183134
rect 471684 182898 472820 183134
rect 473056 182898 473666 183134
rect 473902 182898 482666 183134
rect 482902 182898 491666 183134
rect 491902 182898 500666 183134
rect 500902 182898 509666 183134
rect 509902 182898 511468 183134
rect 511704 182898 512840 183134
rect 513076 182898 513686 183134
rect 513922 182898 522686 183134
rect 522922 182898 531686 183134
rect 531922 182898 540686 183134
rect 540922 182898 549686 183134
rect 549922 182898 551488 183134
rect 551724 182898 552860 183134
rect 553096 182898 553706 183134
rect 553942 182898 562706 183134
rect 562942 182898 571706 183134
rect 571942 182898 573476 183134
rect 573712 182898 578670 183134
rect 578906 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 4582 165454
rect 4818 165218 12232 165454
rect 12468 165218 13038 165454
rect 13274 165218 22038 165454
rect 22274 165218 27588 165454
rect 27824 165218 28240 165454
rect 28476 165218 29046 165454
rect 29282 165218 38046 165454
rect 38282 165218 47046 165454
rect 47282 165218 56046 165454
rect 56282 165218 65046 165454
rect 65282 165218 67608 165454
rect 67844 165218 68260 165454
rect 68496 165218 69066 165454
rect 69302 165218 78066 165454
rect 78302 165218 87066 165454
rect 87302 165218 96066 165454
rect 96302 165218 105066 165454
rect 105302 165218 107628 165454
rect 107864 165218 108280 165454
rect 108516 165218 109086 165454
rect 109322 165218 118086 165454
rect 118322 165218 127086 165454
rect 127322 165218 136086 165454
rect 136322 165218 145086 165454
rect 145322 165218 147648 165454
rect 147884 165218 149300 165454
rect 149536 165218 150106 165454
rect 150342 165218 159106 165454
rect 159342 165218 168106 165454
rect 168342 165218 177106 165454
rect 177342 165218 186106 165454
rect 186342 165218 188668 165454
rect 188904 165218 190320 165454
rect 190556 165218 191126 165454
rect 191362 165218 200126 165454
rect 200362 165218 209126 165454
rect 209362 165218 218126 165454
rect 218362 165218 227126 165454
rect 227362 165218 229688 165454
rect 229924 165218 230340 165454
rect 230576 165218 231146 165454
rect 231382 165218 240146 165454
rect 240382 165218 249146 165454
rect 249382 165218 258146 165454
rect 258382 165218 267146 165454
rect 267382 165218 269708 165454
rect 269944 165218 270360 165454
rect 270596 165218 271166 165454
rect 271402 165218 280166 165454
rect 280402 165218 289166 165454
rect 289402 165218 298166 165454
rect 298402 165218 307166 165454
rect 307402 165218 309728 165454
rect 309964 165218 311380 165454
rect 311616 165218 312186 165454
rect 312422 165218 321186 165454
rect 321422 165218 330186 165454
rect 330422 165218 339186 165454
rect 339422 165218 348186 165454
rect 348422 165218 350748 165454
rect 350984 165218 352400 165454
rect 352636 165218 353206 165454
rect 353442 165218 362206 165454
rect 362442 165218 371206 165454
rect 371442 165218 380206 165454
rect 380442 165218 389206 165454
rect 389442 165218 391768 165454
rect 392004 165218 392420 165454
rect 392656 165218 393226 165454
rect 393462 165218 402226 165454
rect 402462 165218 411226 165454
rect 411462 165218 420226 165454
rect 420462 165218 429226 165454
rect 429462 165218 431788 165454
rect 432024 165218 432440 165454
rect 432676 165218 433246 165454
rect 433482 165218 442246 165454
rect 442482 165218 451246 165454
rect 451482 165218 460246 165454
rect 460482 165218 469246 165454
rect 469482 165218 471808 165454
rect 472044 165218 472460 165454
rect 472696 165218 473266 165454
rect 473502 165218 482266 165454
rect 482502 165218 491266 165454
rect 491502 165218 500266 165454
rect 500502 165218 509266 165454
rect 509502 165218 511828 165454
rect 512064 165218 512480 165454
rect 512716 165218 513286 165454
rect 513522 165218 522286 165454
rect 522522 165218 531286 165454
rect 531522 165218 540286 165454
rect 540522 165218 549286 165454
rect 549522 165218 551848 165454
rect 552084 165218 552500 165454
rect 552736 165218 553306 165454
rect 553542 165218 562306 165454
rect 562542 165218 571306 165454
rect 571542 165218 573836 165454
rect 574072 165218 579470 165454
rect 579706 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 4582 165134
rect 4818 164898 12232 165134
rect 12468 164898 13038 165134
rect 13274 164898 22038 165134
rect 22274 164898 27588 165134
rect 27824 164898 28240 165134
rect 28476 164898 29046 165134
rect 29282 164898 38046 165134
rect 38282 164898 47046 165134
rect 47282 164898 56046 165134
rect 56282 164898 65046 165134
rect 65282 164898 67608 165134
rect 67844 164898 68260 165134
rect 68496 164898 69066 165134
rect 69302 164898 78066 165134
rect 78302 164898 87066 165134
rect 87302 164898 96066 165134
rect 96302 164898 105066 165134
rect 105302 164898 107628 165134
rect 107864 164898 108280 165134
rect 108516 164898 109086 165134
rect 109322 164898 118086 165134
rect 118322 164898 127086 165134
rect 127322 164898 136086 165134
rect 136322 164898 145086 165134
rect 145322 164898 147648 165134
rect 147884 164898 149300 165134
rect 149536 164898 150106 165134
rect 150342 164898 159106 165134
rect 159342 164898 168106 165134
rect 168342 164898 177106 165134
rect 177342 164898 186106 165134
rect 186342 164898 188668 165134
rect 188904 164898 190320 165134
rect 190556 164898 191126 165134
rect 191362 164898 200126 165134
rect 200362 164898 209126 165134
rect 209362 164898 218126 165134
rect 218362 164898 227126 165134
rect 227362 164898 229688 165134
rect 229924 164898 230340 165134
rect 230576 164898 231146 165134
rect 231382 164898 240146 165134
rect 240382 164898 249146 165134
rect 249382 164898 258146 165134
rect 258382 164898 267146 165134
rect 267382 164898 269708 165134
rect 269944 164898 270360 165134
rect 270596 164898 271166 165134
rect 271402 164898 280166 165134
rect 280402 164898 289166 165134
rect 289402 164898 298166 165134
rect 298402 164898 307166 165134
rect 307402 164898 309728 165134
rect 309964 164898 311380 165134
rect 311616 164898 312186 165134
rect 312422 164898 321186 165134
rect 321422 164898 330186 165134
rect 330422 164898 339186 165134
rect 339422 164898 348186 165134
rect 348422 164898 350748 165134
rect 350984 164898 352400 165134
rect 352636 164898 353206 165134
rect 353442 164898 362206 165134
rect 362442 164898 371206 165134
rect 371442 164898 380206 165134
rect 380442 164898 389206 165134
rect 389442 164898 391768 165134
rect 392004 164898 392420 165134
rect 392656 164898 393226 165134
rect 393462 164898 402226 165134
rect 402462 164898 411226 165134
rect 411462 164898 420226 165134
rect 420462 164898 429226 165134
rect 429462 164898 431788 165134
rect 432024 164898 432440 165134
rect 432676 164898 433246 165134
rect 433482 164898 442246 165134
rect 442482 164898 451246 165134
rect 451482 164898 460246 165134
rect 460482 164898 469246 165134
rect 469482 164898 471808 165134
rect 472044 164898 472460 165134
rect 472696 164898 473266 165134
rect 473502 164898 482266 165134
rect 482502 164898 491266 165134
rect 491502 164898 500266 165134
rect 500502 164898 509266 165134
rect 509502 164898 511828 165134
rect 512064 164898 512480 165134
rect 512716 164898 513286 165134
rect 513522 164898 522286 165134
rect 522522 164898 531286 165134
rect 531522 164898 540286 165134
rect 540522 164898 549286 165134
rect 549522 164898 551848 165134
rect 552084 164898 552500 165134
rect 552736 164898 553306 165134
rect 553542 164898 562306 165134
rect 562542 164898 571306 165134
rect 571542 164898 573836 165134
rect 574072 164898 579470 165134
rect 579706 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 5382 147454
rect 5618 147218 12592 147454
rect 12828 147218 13438 147454
rect 13674 147218 22438 147454
rect 22674 147218 27228 147454
rect 27464 147218 28600 147454
rect 28836 147218 29446 147454
rect 29682 147218 38446 147454
rect 38682 147218 47446 147454
rect 47682 147218 56446 147454
rect 56682 147218 65446 147454
rect 65682 147218 67248 147454
rect 67484 147218 68620 147454
rect 68856 147218 69466 147454
rect 69702 147218 78466 147454
rect 78702 147218 87466 147454
rect 87702 147218 96466 147454
rect 96702 147218 105466 147454
rect 105702 147218 107268 147454
rect 107504 147218 108640 147454
rect 108876 147218 109486 147454
rect 109722 147218 118486 147454
rect 118722 147218 127486 147454
rect 127722 147218 136486 147454
rect 136722 147218 145486 147454
rect 145722 147218 147288 147454
rect 147524 147218 149660 147454
rect 149896 147218 150506 147454
rect 150742 147218 159506 147454
rect 159742 147218 168506 147454
rect 168742 147218 177506 147454
rect 177742 147218 186506 147454
rect 186742 147218 188308 147454
rect 188544 147218 190680 147454
rect 190916 147218 191526 147454
rect 191762 147218 200526 147454
rect 200762 147218 209526 147454
rect 209762 147218 218526 147454
rect 218762 147218 227526 147454
rect 227762 147218 229328 147454
rect 229564 147218 230700 147454
rect 230936 147218 231546 147454
rect 231782 147218 240546 147454
rect 240782 147218 249546 147454
rect 249782 147218 258546 147454
rect 258782 147218 267546 147454
rect 267782 147218 269348 147454
rect 269584 147218 270720 147454
rect 270956 147218 271566 147454
rect 271802 147218 280566 147454
rect 280802 147218 289566 147454
rect 289802 147218 298566 147454
rect 298802 147218 307566 147454
rect 307802 147218 309368 147454
rect 309604 147218 311740 147454
rect 311976 147218 312586 147454
rect 312822 147218 321586 147454
rect 321822 147218 330586 147454
rect 330822 147218 339586 147454
rect 339822 147218 348586 147454
rect 348822 147218 350388 147454
rect 350624 147218 352760 147454
rect 352996 147218 353606 147454
rect 353842 147218 362606 147454
rect 362842 147218 371606 147454
rect 371842 147218 380606 147454
rect 380842 147218 389606 147454
rect 389842 147218 391408 147454
rect 391644 147218 392780 147454
rect 393016 147218 393626 147454
rect 393862 147218 402626 147454
rect 402862 147218 411626 147454
rect 411862 147218 420626 147454
rect 420862 147218 429626 147454
rect 429862 147218 431428 147454
rect 431664 147218 432800 147454
rect 433036 147218 433646 147454
rect 433882 147218 442646 147454
rect 442882 147218 451646 147454
rect 451882 147218 460646 147454
rect 460882 147218 469646 147454
rect 469882 147218 471448 147454
rect 471684 147218 472820 147454
rect 473056 147218 473666 147454
rect 473902 147218 482666 147454
rect 482902 147218 491666 147454
rect 491902 147218 500666 147454
rect 500902 147218 509666 147454
rect 509902 147218 511468 147454
rect 511704 147218 512840 147454
rect 513076 147218 513686 147454
rect 513922 147218 522686 147454
rect 522922 147218 531686 147454
rect 531922 147218 540686 147454
rect 540922 147218 549686 147454
rect 549922 147218 551488 147454
rect 551724 147218 552860 147454
rect 553096 147218 553706 147454
rect 553942 147218 562706 147454
rect 562942 147218 571706 147454
rect 571942 147218 573476 147454
rect 573712 147218 578670 147454
rect 578906 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 5382 147134
rect 5618 146898 12592 147134
rect 12828 146898 13438 147134
rect 13674 146898 22438 147134
rect 22674 146898 27228 147134
rect 27464 146898 28600 147134
rect 28836 146898 29446 147134
rect 29682 146898 38446 147134
rect 38682 146898 47446 147134
rect 47682 146898 56446 147134
rect 56682 146898 65446 147134
rect 65682 146898 67248 147134
rect 67484 146898 68620 147134
rect 68856 146898 69466 147134
rect 69702 146898 78466 147134
rect 78702 146898 87466 147134
rect 87702 146898 96466 147134
rect 96702 146898 105466 147134
rect 105702 146898 107268 147134
rect 107504 146898 108640 147134
rect 108876 146898 109486 147134
rect 109722 146898 118486 147134
rect 118722 146898 127486 147134
rect 127722 146898 136486 147134
rect 136722 146898 145486 147134
rect 145722 146898 147288 147134
rect 147524 146898 149660 147134
rect 149896 146898 150506 147134
rect 150742 146898 159506 147134
rect 159742 146898 168506 147134
rect 168742 146898 177506 147134
rect 177742 146898 186506 147134
rect 186742 146898 188308 147134
rect 188544 146898 190680 147134
rect 190916 146898 191526 147134
rect 191762 146898 200526 147134
rect 200762 146898 209526 147134
rect 209762 146898 218526 147134
rect 218762 146898 227526 147134
rect 227762 146898 229328 147134
rect 229564 146898 230700 147134
rect 230936 146898 231546 147134
rect 231782 146898 240546 147134
rect 240782 146898 249546 147134
rect 249782 146898 258546 147134
rect 258782 146898 267546 147134
rect 267782 146898 269348 147134
rect 269584 146898 270720 147134
rect 270956 146898 271566 147134
rect 271802 146898 280566 147134
rect 280802 146898 289566 147134
rect 289802 146898 298566 147134
rect 298802 146898 307566 147134
rect 307802 146898 309368 147134
rect 309604 146898 311740 147134
rect 311976 146898 312586 147134
rect 312822 146898 321586 147134
rect 321822 146898 330586 147134
rect 330822 146898 339586 147134
rect 339822 146898 348586 147134
rect 348822 146898 350388 147134
rect 350624 146898 352760 147134
rect 352996 146898 353606 147134
rect 353842 146898 362606 147134
rect 362842 146898 371606 147134
rect 371842 146898 380606 147134
rect 380842 146898 389606 147134
rect 389842 146898 391408 147134
rect 391644 146898 392780 147134
rect 393016 146898 393626 147134
rect 393862 146898 402626 147134
rect 402862 146898 411626 147134
rect 411862 146898 420626 147134
rect 420862 146898 429626 147134
rect 429862 146898 431428 147134
rect 431664 146898 432800 147134
rect 433036 146898 433646 147134
rect 433882 146898 442646 147134
rect 442882 146898 451646 147134
rect 451882 146898 460646 147134
rect 460882 146898 469646 147134
rect 469882 146898 471448 147134
rect 471684 146898 472820 147134
rect 473056 146898 473666 147134
rect 473902 146898 482666 147134
rect 482902 146898 491666 147134
rect 491902 146898 500666 147134
rect 500902 146898 509666 147134
rect 509902 146898 511468 147134
rect 511704 146898 512840 147134
rect 513076 146898 513686 147134
rect 513922 146898 522686 147134
rect 522922 146898 531686 147134
rect 531922 146898 540686 147134
rect 540922 146898 549686 147134
rect 549922 146898 551488 147134
rect 551724 146898 552860 147134
rect 553096 146898 553706 147134
rect 553942 146898 562706 147134
rect 562942 146898 571706 147134
rect 571942 146898 573476 147134
rect 573712 146898 578670 147134
rect 578906 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 4582 129454
rect 4818 129218 12232 129454
rect 12468 129218 13038 129454
rect 13274 129218 22038 129454
rect 22274 129218 27588 129454
rect 27824 129218 28240 129454
rect 28476 129218 29046 129454
rect 29282 129218 38046 129454
rect 38282 129218 47046 129454
rect 47282 129218 56046 129454
rect 56282 129218 65046 129454
rect 65282 129218 67608 129454
rect 67844 129218 68260 129454
rect 68496 129218 69066 129454
rect 69302 129218 78066 129454
rect 78302 129218 87066 129454
rect 87302 129218 96066 129454
rect 96302 129218 105066 129454
rect 105302 129218 107628 129454
rect 107864 129218 108280 129454
rect 108516 129218 109086 129454
rect 109322 129218 118086 129454
rect 118322 129218 127086 129454
rect 127322 129218 136086 129454
rect 136322 129218 145086 129454
rect 145322 129218 147648 129454
rect 147884 129218 149300 129454
rect 149536 129218 150106 129454
rect 150342 129218 159106 129454
rect 159342 129218 168106 129454
rect 168342 129218 177106 129454
rect 177342 129218 186106 129454
rect 186342 129218 188668 129454
rect 188904 129218 190320 129454
rect 190556 129218 191126 129454
rect 191362 129218 200126 129454
rect 200362 129218 209126 129454
rect 209362 129218 218126 129454
rect 218362 129218 227126 129454
rect 227362 129218 229688 129454
rect 229924 129218 230340 129454
rect 230576 129218 231146 129454
rect 231382 129218 240146 129454
rect 240382 129218 249146 129454
rect 249382 129218 258146 129454
rect 258382 129218 267146 129454
rect 267382 129218 269708 129454
rect 269944 129218 270360 129454
rect 270596 129218 271166 129454
rect 271402 129218 280166 129454
rect 280402 129218 289166 129454
rect 289402 129218 298166 129454
rect 298402 129218 307166 129454
rect 307402 129218 309728 129454
rect 309964 129218 311380 129454
rect 311616 129218 312186 129454
rect 312422 129218 321186 129454
rect 321422 129218 330186 129454
rect 330422 129218 339186 129454
rect 339422 129218 348186 129454
rect 348422 129218 350748 129454
rect 350984 129218 352400 129454
rect 352636 129218 353206 129454
rect 353442 129218 362206 129454
rect 362442 129218 371206 129454
rect 371442 129218 380206 129454
rect 380442 129218 389206 129454
rect 389442 129218 391768 129454
rect 392004 129218 392420 129454
rect 392656 129218 393226 129454
rect 393462 129218 402226 129454
rect 402462 129218 411226 129454
rect 411462 129218 420226 129454
rect 420462 129218 429226 129454
rect 429462 129218 431788 129454
rect 432024 129218 432440 129454
rect 432676 129218 433246 129454
rect 433482 129218 442246 129454
rect 442482 129218 451246 129454
rect 451482 129218 460246 129454
rect 460482 129218 469246 129454
rect 469482 129218 471808 129454
rect 472044 129218 472460 129454
rect 472696 129218 473266 129454
rect 473502 129218 482266 129454
rect 482502 129218 491266 129454
rect 491502 129218 500266 129454
rect 500502 129218 509266 129454
rect 509502 129218 511828 129454
rect 512064 129218 512480 129454
rect 512716 129218 513286 129454
rect 513522 129218 522286 129454
rect 522522 129218 531286 129454
rect 531522 129218 540286 129454
rect 540522 129218 549286 129454
rect 549522 129218 551848 129454
rect 552084 129218 552500 129454
rect 552736 129218 553306 129454
rect 553542 129218 562306 129454
rect 562542 129218 571306 129454
rect 571542 129218 573836 129454
rect 574072 129218 579470 129454
rect 579706 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 4582 129134
rect 4818 128898 12232 129134
rect 12468 128898 13038 129134
rect 13274 128898 22038 129134
rect 22274 128898 27588 129134
rect 27824 128898 28240 129134
rect 28476 128898 29046 129134
rect 29282 128898 38046 129134
rect 38282 128898 47046 129134
rect 47282 128898 56046 129134
rect 56282 128898 65046 129134
rect 65282 128898 67608 129134
rect 67844 128898 68260 129134
rect 68496 128898 69066 129134
rect 69302 128898 78066 129134
rect 78302 128898 87066 129134
rect 87302 128898 96066 129134
rect 96302 128898 105066 129134
rect 105302 128898 107628 129134
rect 107864 128898 108280 129134
rect 108516 128898 109086 129134
rect 109322 128898 118086 129134
rect 118322 128898 127086 129134
rect 127322 128898 136086 129134
rect 136322 128898 145086 129134
rect 145322 128898 147648 129134
rect 147884 128898 149300 129134
rect 149536 128898 150106 129134
rect 150342 128898 159106 129134
rect 159342 128898 168106 129134
rect 168342 128898 177106 129134
rect 177342 128898 186106 129134
rect 186342 128898 188668 129134
rect 188904 128898 190320 129134
rect 190556 128898 191126 129134
rect 191362 128898 200126 129134
rect 200362 128898 209126 129134
rect 209362 128898 218126 129134
rect 218362 128898 227126 129134
rect 227362 128898 229688 129134
rect 229924 128898 230340 129134
rect 230576 128898 231146 129134
rect 231382 128898 240146 129134
rect 240382 128898 249146 129134
rect 249382 128898 258146 129134
rect 258382 128898 267146 129134
rect 267382 128898 269708 129134
rect 269944 128898 270360 129134
rect 270596 128898 271166 129134
rect 271402 128898 280166 129134
rect 280402 128898 289166 129134
rect 289402 128898 298166 129134
rect 298402 128898 307166 129134
rect 307402 128898 309728 129134
rect 309964 128898 311380 129134
rect 311616 128898 312186 129134
rect 312422 128898 321186 129134
rect 321422 128898 330186 129134
rect 330422 128898 339186 129134
rect 339422 128898 348186 129134
rect 348422 128898 350748 129134
rect 350984 128898 352400 129134
rect 352636 128898 353206 129134
rect 353442 128898 362206 129134
rect 362442 128898 371206 129134
rect 371442 128898 380206 129134
rect 380442 128898 389206 129134
rect 389442 128898 391768 129134
rect 392004 128898 392420 129134
rect 392656 128898 393226 129134
rect 393462 128898 402226 129134
rect 402462 128898 411226 129134
rect 411462 128898 420226 129134
rect 420462 128898 429226 129134
rect 429462 128898 431788 129134
rect 432024 128898 432440 129134
rect 432676 128898 433246 129134
rect 433482 128898 442246 129134
rect 442482 128898 451246 129134
rect 451482 128898 460246 129134
rect 460482 128898 469246 129134
rect 469482 128898 471808 129134
rect 472044 128898 472460 129134
rect 472696 128898 473266 129134
rect 473502 128898 482266 129134
rect 482502 128898 491266 129134
rect 491502 128898 500266 129134
rect 500502 128898 509266 129134
rect 509502 128898 511828 129134
rect 512064 128898 512480 129134
rect 512716 128898 513286 129134
rect 513522 128898 522286 129134
rect 522522 128898 531286 129134
rect 531522 128898 540286 129134
rect 540522 128898 549286 129134
rect 549522 128898 551848 129134
rect 552084 128898 552500 129134
rect 552736 128898 553306 129134
rect 553542 128898 562306 129134
rect 562542 128898 571306 129134
rect 571542 128898 573836 129134
rect 574072 128898 579470 129134
rect 579706 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 5382 111454
rect 5618 111218 12592 111454
rect 12828 111218 13438 111454
rect 13674 111218 22438 111454
rect 22674 111218 27228 111454
rect 27464 111218 28600 111454
rect 28836 111218 29446 111454
rect 29682 111218 38446 111454
rect 38682 111218 47446 111454
rect 47682 111218 56446 111454
rect 56682 111218 65446 111454
rect 65682 111218 67248 111454
rect 67484 111218 68620 111454
rect 68856 111218 69466 111454
rect 69702 111218 78466 111454
rect 78702 111218 87466 111454
rect 87702 111218 96466 111454
rect 96702 111218 105466 111454
rect 105702 111218 107268 111454
rect 107504 111218 108640 111454
rect 108876 111218 109486 111454
rect 109722 111218 118486 111454
rect 118722 111218 127486 111454
rect 127722 111218 136486 111454
rect 136722 111218 145486 111454
rect 145722 111218 147288 111454
rect 147524 111218 149660 111454
rect 149896 111218 150506 111454
rect 150742 111218 159506 111454
rect 159742 111218 168506 111454
rect 168742 111218 177506 111454
rect 177742 111218 186506 111454
rect 186742 111218 188308 111454
rect 188544 111218 190680 111454
rect 190916 111218 191526 111454
rect 191762 111218 200526 111454
rect 200762 111218 209526 111454
rect 209762 111218 218526 111454
rect 218762 111218 227526 111454
rect 227762 111218 229328 111454
rect 229564 111218 230700 111454
rect 230936 111218 231546 111454
rect 231782 111218 240546 111454
rect 240782 111218 249546 111454
rect 249782 111218 258546 111454
rect 258782 111218 267546 111454
rect 267782 111218 269348 111454
rect 269584 111218 270720 111454
rect 270956 111218 271566 111454
rect 271802 111218 280566 111454
rect 280802 111218 289566 111454
rect 289802 111218 298566 111454
rect 298802 111218 307566 111454
rect 307802 111218 309368 111454
rect 309604 111218 311740 111454
rect 311976 111218 312586 111454
rect 312822 111218 321586 111454
rect 321822 111218 330586 111454
rect 330822 111218 339586 111454
rect 339822 111218 348586 111454
rect 348822 111218 350388 111454
rect 350624 111218 352760 111454
rect 352996 111218 353606 111454
rect 353842 111218 362606 111454
rect 362842 111218 371606 111454
rect 371842 111218 380606 111454
rect 380842 111218 389606 111454
rect 389842 111218 391408 111454
rect 391644 111218 392780 111454
rect 393016 111218 393626 111454
rect 393862 111218 402626 111454
rect 402862 111218 411626 111454
rect 411862 111218 420626 111454
rect 420862 111218 429626 111454
rect 429862 111218 431428 111454
rect 431664 111218 432800 111454
rect 433036 111218 433646 111454
rect 433882 111218 442646 111454
rect 442882 111218 451646 111454
rect 451882 111218 460646 111454
rect 460882 111218 469646 111454
rect 469882 111218 471448 111454
rect 471684 111218 472820 111454
rect 473056 111218 473666 111454
rect 473902 111218 482666 111454
rect 482902 111218 491666 111454
rect 491902 111218 500666 111454
rect 500902 111218 509666 111454
rect 509902 111218 511468 111454
rect 511704 111218 512840 111454
rect 513076 111218 513686 111454
rect 513922 111218 522686 111454
rect 522922 111218 531686 111454
rect 531922 111218 540686 111454
rect 540922 111218 549686 111454
rect 549922 111218 551488 111454
rect 551724 111218 552860 111454
rect 553096 111218 553706 111454
rect 553942 111218 562706 111454
rect 562942 111218 571706 111454
rect 571942 111218 573476 111454
rect 573712 111218 578670 111454
rect 578906 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 5382 111134
rect 5618 110898 12592 111134
rect 12828 110898 13438 111134
rect 13674 110898 22438 111134
rect 22674 110898 27228 111134
rect 27464 110898 28600 111134
rect 28836 110898 29446 111134
rect 29682 110898 38446 111134
rect 38682 110898 47446 111134
rect 47682 110898 56446 111134
rect 56682 110898 65446 111134
rect 65682 110898 67248 111134
rect 67484 110898 68620 111134
rect 68856 110898 69466 111134
rect 69702 110898 78466 111134
rect 78702 110898 87466 111134
rect 87702 110898 96466 111134
rect 96702 110898 105466 111134
rect 105702 110898 107268 111134
rect 107504 110898 108640 111134
rect 108876 110898 109486 111134
rect 109722 110898 118486 111134
rect 118722 110898 127486 111134
rect 127722 110898 136486 111134
rect 136722 110898 145486 111134
rect 145722 110898 147288 111134
rect 147524 110898 149660 111134
rect 149896 110898 150506 111134
rect 150742 110898 159506 111134
rect 159742 110898 168506 111134
rect 168742 110898 177506 111134
rect 177742 110898 186506 111134
rect 186742 110898 188308 111134
rect 188544 110898 190680 111134
rect 190916 110898 191526 111134
rect 191762 110898 200526 111134
rect 200762 110898 209526 111134
rect 209762 110898 218526 111134
rect 218762 110898 227526 111134
rect 227762 110898 229328 111134
rect 229564 110898 230700 111134
rect 230936 110898 231546 111134
rect 231782 110898 240546 111134
rect 240782 110898 249546 111134
rect 249782 110898 258546 111134
rect 258782 110898 267546 111134
rect 267782 110898 269348 111134
rect 269584 110898 270720 111134
rect 270956 110898 271566 111134
rect 271802 110898 280566 111134
rect 280802 110898 289566 111134
rect 289802 110898 298566 111134
rect 298802 110898 307566 111134
rect 307802 110898 309368 111134
rect 309604 110898 311740 111134
rect 311976 110898 312586 111134
rect 312822 110898 321586 111134
rect 321822 110898 330586 111134
rect 330822 110898 339586 111134
rect 339822 110898 348586 111134
rect 348822 110898 350388 111134
rect 350624 110898 352760 111134
rect 352996 110898 353606 111134
rect 353842 110898 362606 111134
rect 362842 110898 371606 111134
rect 371842 110898 380606 111134
rect 380842 110898 389606 111134
rect 389842 110898 391408 111134
rect 391644 110898 392780 111134
rect 393016 110898 393626 111134
rect 393862 110898 402626 111134
rect 402862 110898 411626 111134
rect 411862 110898 420626 111134
rect 420862 110898 429626 111134
rect 429862 110898 431428 111134
rect 431664 110898 432800 111134
rect 433036 110898 433646 111134
rect 433882 110898 442646 111134
rect 442882 110898 451646 111134
rect 451882 110898 460646 111134
rect 460882 110898 469646 111134
rect 469882 110898 471448 111134
rect 471684 110898 472820 111134
rect 473056 110898 473666 111134
rect 473902 110898 482666 111134
rect 482902 110898 491666 111134
rect 491902 110898 500666 111134
rect 500902 110898 509666 111134
rect 509902 110898 511468 111134
rect 511704 110898 512840 111134
rect 513076 110898 513686 111134
rect 513922 110898 522686 111134
rect 522922 110898 531686 111134
rect 531922 110898 540686 111134
rect 540922 110898 549686 111134
rect 549922 110898 551488 111134
rect 551724 110898 552860 111134
rect 553096 110898 553706 111134
rect 553942 110898 562706 111134
rect 562942 110898 571706 111134
rect 571942 110898 573476 111134
rect 573712 110898 578670 111134
rect 578906 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 4582 93454
rect 4818 93218 12232 93454
rect 12468 93218 13038 93454
rect 13274 93218 22038 93454
rect 22274 93218 27588 93454
rect 27824 93218 28240 93454
rect 28476 93218 29046 93454
rect 29282 93218 38046 93454
rect 38282 93218 47046 93454
rect 47282 93218 56046 93454
rect 56282 93218 65046 93454
rect 65282 93218 67608 93454
rect 67844 93218 68260 93454
rect 68496 93218 69066 93454
rect 69302 93218 78066 93454
rect 78302 93218 87066 93454
rect 87302 93218 96066 93454
rect 96302 93218 105066 93454
rect 105302 93218 107628 93454
rect 107864 93218 108280 93454
rect 108516 93218 109086 93454
rect 109322 93218 118086 93454
rect 118322 93218 127086 93454
rect 127322 93218 136086 93454
rect 136322 93218 145086 93454
rect 145322 93218 147648 93454
rect 147884 93218 149300 93454
rect 149536 93218 150106 93454
rect 150342 93218 159106 93454
rect 159342 93218 168106 93454
rect 168342 93218 177106 93454
rect 177342 93218 186106 93454
rect 186342 93218 188668 93454
rect 188904 93218 190320 93454
rect 190556 93218 191126 93454
rect 191362 93218 200126 93454
rect 200362 93218 209126 93454
rect 209362 93218 218126 93454
rect 218362 93218 227126 93454
rect 227362 93218 229688 93454
rect 229924 93218 230340 93454
rect 230576 93218 231146 93454
rect 231382 93218 240146 93454
rect 240382 93218 249146 93454
rect 249382 93218 258146 93454
rect 258382 93218 267146 93454
rect 267382 93218 269708 93454
rect 269944 93218 270360 93454
rect 270596 93218 271166 93454
rect 271402 93218 280166 93454
rect 280402 93218 289166 93454
rect 289402 93218 298166 93454
rect 298402 93218 307166 93454
rect 307402 93218 309728 93454
rect 309964 93218 311380 93454
rect 311616 93218 312186 93454
rect 312422 93218 321186 93454
rect 321422 93218 330186 93454
rect 330422 93218 339186 93454
rect 339422 93218 348186 93454
rect 348422 93218 350748 93454
rect 350984 93218 352400 93454
rect 352636 93218 353206 93454
rect 353442 93218 362206 93454
rect 362442 93218 371206 93454
rect 371442 93218 380206 93454
rect 380442 93218 389206 93454
rect 389442 93218 391768 93454
rect 392004 93218 392420 93454
rect 392656 93218 393226 93454
rect 393462 93218 402226 93454
rect 402462 93218 411226 93454
rect 411462 93218 420226 93454
rect 420462 93218 429226 93454
rect 429462 93218 431788 93454
rect 432024 93218 432440 93454
rect 432676 93218 433246 93454
rect 433482 93218 442246 93454
rect 442482 93218 451246 93454
rect 451482 93218 460246 93454
rect 460482 93218 469246 93454
rect 469482 93218 471808 93454
rect 472044 93218 472460 93454
rect 472696 93218 473266 93454
rect 473502 93218 482266 93454
rect 482502 93218 491266 93454
rect 491502 93218 500266 93454
rect 500502 93218 509266 93454
rect 509502 93218 511828 93454
rect 512064 93218 512480 93454
rect 512716 93218 513286 93454
rect 513522 93218 522286 93454
rect 522522 93218 531286 93454
rect 531522 93218 540286 93454
rect 540522 93218 549286 93454
rect 549522 93218 551848 93454
rect 552084 93218 552500 93454
rect 552736 93218 553306 93454
rect 553542 93218 562306 93454
rect 562542 93218 571306 93454
rect 571542 93218 573836 93454
rect 574072 93218 579470 93454
rect 579706 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 4582 93134
rect 4818 92898 12232 93134
rect 12468 92898 13038 93134
rect 13274 92898 22038 93134
rect 22274 92898 27588 93134
rect 27824 92898 28240 93134
rect 28476 92898 29046 93134
rect 29282 92898 38046 93134
rect 38282 92898 47046 93134
rect 47282 92898 56046 93134
rect 56282 92898 65046 93134
rect 65282 92898 67608 93134
rect 67844 92898 68260 93134
rect 68496 92898 69066 93134
rect 69302 92898 78066 93134
rect 78302 92898 87066 93134
rect 87302 92898 96066 93134
rect 96302 92898 105066 93134
rect 105302 92898 107628 93134
rect 107864 92898 108280 93134
rect 108516 92898 109086 93134
rect 109322 92898 118086 93134
rect 118322 92898 127086 93134
rect 127322 92898 136086 93134
rect 136322 92898 145086 93134
rect 145322 92898 147648 93134
rect 147884 92898 149300 93134
rect 149536 92898 150106 93134
rect 150342 92898 159106 93134
rect 159342 92898 168106 93134
rect 168342 92898 177106 93134
rect 177342 92898 186106 93134
rect 186342 92898 188668 93134
rect 188904 92898 190320 93134
rect 190556 92898 191126 93134
rect 191362 92898 200126 93134
rect 200362 92898 209126 93134
rect 209362 92898 218126 93134
rect 218362 92898 227126 93134
rect 227362 92898 229688 93134
rect 229924 92898 230340 93134
rect 230576 92898 231146 93134
rect 231382 92898 240146 93134
rect 240382 92898 249146 93134
rect 249382 92898 258146 93134
rect 258382 92898 267146 93134
rect 267382 92898 269708 93134
rect 269944 92898 270360 93134
rect 270596 92898 271166 93134
rect 271402 92898 280166 93134
rect 280402 92898 289166 93134
rect 289402 92898 298166 93134
rect 298402 92898 307166 93134
rect 307402 92898 309728 93134
rect 309964 92898 311380 93134
rect 311616 92898 312186 93134
rect 312422 92898 321186 93134
rect 321422 92898 330186 93134
rect 330422 92898 339186 93134
rect 339422 92898 348186 93134
rect 348422 92898 350748 93134
rect 350984 92898 352400 93134
rect 352636 92898 353206 93134
rect 353442 92898 362206 93134
rect 362442 92898 371206 93134
rect 371442 92898 380206 93134
rect 380442 92898 389206 93134
rect 389442 92898 391768 93134
rect 392004 92898 392420 93134
rect 392656 92898 393226 93134
rect 393462 92898 402226 93134
rect 402462 92898 411226 93134
rect 411462 92898 420226 93134
rect 420462 92898 429226 93134
rect 429462 92898 431788 93134
rect 432024 92898 432440 93134
rect 432676 92898 433246 93134
rect 433482 92898 442246 93134
rect 442482 92898 451246 93134
rect 451482 92898 460246 93134
rect 460482 92898 469246 93134
rect 469482 92898 471808 93134
rect 472044 92898 472460 93134
rect 472696 92898 473266 93134
rect 473502 92898 482266 93134
rect 482502 92898 491266 93134
rect 491502 92898 500266 93134
rect 500502 92898 509266 93134
rect 509502 92898 511828 93134
rect 512064 92898 512480 93134
rect 512716 92898 513286 93134
rect 513522 92898 522286 93134
rect 522522 92898 531286 93134
rect 531522 92898 540286 93134
rect 540522 92898 549286 93134
rect 549522 92898 551848 93134
rect 552084 92898 552500 93134
rect 552736 92898 553306 93134
rect 553542 92898 562306 93134
rect 562542 92898 571306 93134
rect 571542 92898 573836 93134
rect 574072 92898 579470 93134
rect 579706 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 5382 75454
rect 5618 75218 12592 75454
rect 12828 75218 13438 75454
rect 13674 75218 22438 75454
rect 22674 75218 27228 75454
rect 27464 75218 28600 75454
rect 28836 75218 29446 75454
rect 29682 75218 38446 75454
rect 38682 75218 47446 75454
rect 47682 75218 56446 75454
rect 56682 75218 65446 75454
rect 65682 75218 67248 75454
rect 67484 75218 68620 75454
rect 68856 75218 69466 75454
rect 69702 75218 78466 75454
rect 78702 75218 87466 75454
rect 87702 75218 96466 75454
rect 96702 75218 105466 75454
rect 105702 75218 107268 75454
rect 107504 75218 108640 75454
rect 108876 75218 109486 75454
rect 109722 75218 118486 75454
rect 118722 75218 127486 75454
rect 127722 75218 136486 75454
rect 136722 75218 145486 75454
rect 145722 75218 147288 75454
rect 147524 75218 149660 75454
rect 149896 75218 150506 75454
rect 150742 75218 159506 75454
rect 159742 75218 168506 75454
rect 168742 75218 177506 75454
rect 177742 75218 186506 75454
rect 186742 75218 188308 75454
rect 188544 75218 190680 75454
rect 190916 75218 191526 75454
rect 191762 75218 200526 75454
rect 200762 75218 209526 75454
rect 209762 75218 218526 75454
rect 218762 75218 227526 75454
rect 227762 75218 229328 75454
rect 229564 75218 230700 75454
rect 230936 75218 231546 75454
rect 231782 75218 240546 75454
rect 240782 75218 249546 75454
rect 249782 75218 258546 75454
rect 258782 75218 267546 75454
rect 267782 75218 269348 75454
rect 269584 75218 270720 75454
rect 270956 75218 271566 75454
rect 271802 75218 280566 75454
rect 280802 75218 289566 75454
rect 289802 75218 298566 75454
rect 298802 75218 307566 75454
rect 307802 75218 309368 75454
rect 309604 75218 311740 75454
rect 311976 75218 312586 75454
rect 312822 75218 321586 75454
rect 321822 75218 330586 75454
rect 330822 75218 339586 75454
rect 339822 75218 348586 75454
rect 348822 75218 350388 75454
rect 350624 75218 352760 75454
rect 352996 75218 353606 75454
rect 353842 75218 362606 75454
rect 362842 75218 371606 75454
rect 371842 75218 380606 75454
rect 380842 75218 389606 75454
rect 389842 75218 391408 75454
rect 391644 75218 392780 75454
rect 393016 75218 393626 75454
rect 393862 75218 402626 75454
rect 402862 75218 411626 75454
rect 411862 75218 420626 75454
rect 420862 75218 429626 75454
rect 429862 75218 431428 75454
rect 431664 75218 432800 75454
rect 433036 75218 433646 75454
rect 433882 75218 442646 75454
rect 442882 75218 451646 75454
rect 451882 75218 460646 75454
rect 460882 75218 469646 75454
rect 469882 75218 471448 75454
rect 471684 75218 472820 75454
rect 473056 75218 473666 75454
rect 473902 75218 482666 75454
rect 482902 75218 491666 75454
rect 491902 75218 500666 75454
rect 500902 75218 509666 75454
rect 509902 75218 511468 75454
rect 511704 75218 512840 75454
rect 513076 75218 513686 75454
rect 513922 75218 522686 75454
rect 522922 75218 531686 75454
rect 531922 75218 540686 75454
rect 540922 75218 549686 75454
rect 549922 75218 551488 75454
rect 551724 75218 552860 75454
rect 553096 75218 553706 75454
rect 553942 75218 562706 75454
rect 562942 75218 571706 75454
rect 571942 75218 573476 75454
rect 573712 75218 578670 75454
rect 578906 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 5382 75134
rect 5618 74898 12592 75134
rect 12828 74898 13438 75134
rect 13674 74898 22438 75134
rect 22674 74898 27228 75134
rect 27464 74898 28600 75134
rect 28836 74898 29446 75134
rect 29682 74898 38446 75134
rect 38682 74898 47446 75134
rect 47682 74898 56446 75134
rect 56682 74898 65446 75134
rect 65682 74898 67248 75134
rect 67484 74898 68620 75134
rect 68856 74898 69466 75134
rect 69702 74898 78466 75134
rect 78702 74898 87466 75134
rect 87702 74898 96466 75134
rect 96702 74898 105466 75134
rect 105702 74898 107268 75134
rect 107504 74898 108640 75134
rect 108876 74898 109486 75134
rect 109722 74898 118486 75134
rect 118722 74898 127486 75134
rect 127722 74898 136486 75134
rect 136722 74898 145486 75134
rect 145722 74898 147288 75134
rect 147524 74898 149660 75134
rect 149896 74898 150506 75134
rect 150742 74898 159506 75134
rect 159742 74898 168506 75134
rect 168742 74898 177506 75134
rect 177742 74898 186506 75134
rect 186742 74898 188308 75134
rect 188544 74898 190680 75134
rect 190916 74898 191526 75134
rect 191762 74898 200526 75134
rect 200762 74898 209526 75134
rect 209762 74898 218526 75134
rect 218762 74898 227526 75134
rect 227762 74898 229328 75134
rect 229564 74898 230700 75134
rect 230936 74898 231546 75134
rect 231782 74898 240546 75134
rect 240782 74898 249546 75134
rect 249782 74898 258546 75134
rect 258782 74898 267546 75134
rect 267782 74898 269348 75134
rect 269584 74898 270720 75134
rect 270956 74898 271566 75134
rect 271802 74898 280566 75134
rect 280802 74898 289566 75134
rect 289802 74898 298566 75134
rect 298802 74898 307566 75134
rect 307802 74898 309368 75134
rect 309604 74898 311740 75134
rect 311976 74898 312586 75134
rect 312822 74898 321586 75134
rect 321822 74898 330586 75134
rect 330822 74898 339586 75134
rect 339822 74898 348586 75134
rect 348822 74898 350388 75134
rect 350624 74898 352760 75134
rect 352996 74898 353606 75134
rect 353842 74898 362606 75134
rect 362842 74898 371606 75134
rect 371842 74898 380606 75134
rect 380842 74898 389606 75134
rect 389842 74898 391408 75134
rect 391644 74898 392780 75134
rect 393016 74898 393626 75134
rect 393862 74898 402626 75134
rect 402862 74898 411626 75134
rect 411862 74898 420626 75134
rect 420862 74898 429626 75134
rect 429862 74898 431428 75134
rect 431664 74898 432800 75134
rect 433036 74898 433646 75134
rect 433882 74898 442646 75134
rect 442882 74898 451646 75134
rect 451882 74898 460646 75134
rect 460882 74898 469646 75134
rect 469882 74898 471448 75134
rect 471684 74898 472820 75134
rect 473056 74898 473666 75134
rect 473902 74898 482666 75134
rect 482902 74898 491666 75134
rect 491902 74898 500666 75134
rect 500902 74898 509666 75134
rect 509902 74898 511468 75134
rect 511704 74898 512840 75134
rect 513076 74898 513686 75134
rect 513922 74898 522686 75134
rect 522922 74898 531686 75134
rect 531922 74898 540686 75134
rect 540922 74898 549686 75134
rect 549922 74898 551488 75134
rect 551724 74898 552860 75134
rect 553096 74898 553706 75134
rect 553942 74898 562706 75134
rect 562942 74898 571706 75134
rect 571942 74898 573476 75134
rect 573712 74898 578670 75134
rect 578906 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 4582 57454
rect 4818 57218 28240 57454
rect 28476 57218 29046 57454
rect 29282 57218 38046 57454
rect 38282 57218 47046 57454
rect 47282 57218 56046 57454
rect 56282 57218 65046 57454
rect 65282 57218 67608 57454
rect 67844 57218 68260 57454
rect 68496 57218 69066 57454
rect 69302 57218 78066 57454
rect 78302 57218 87066 57454
rect 87302 57218 96066 57454
rect 96302 57218 105066 57454
rect 105302 57218 107628 57454
rect 107864 57218 108280 57454
rect 108516 57218 109086 57454
rect 109322 57218 118086 57454
rect 118322 57218 127086 57454
rect 127322 57218 136086 57454
rect 136322 57218 145086 57454
rect 145322 57218 147648 57454
rect 147884 57218 149300 57454
rect 149536 57218 150106 57454
rect 150342 57218 159106 57454
rect 159342 57218 168106 57454
rect 168342 57218 177106 57454
rect 177342 57218 186106 57454
rect 186342 57218 188668 57454
rect 188904 57218 190320 57454
rect 190556 57218 191126 57454
rect 191362 57218 200126 57454
rect 200362 57218 209126 57454
rect 209362 57218 218126 57454
rect 218362 57218 227126 57454
rect 227362 57218 229688 57454
rect 229924 57218 230340 57454
rect 230576 57218 231146 57454
rect 231382 57218 240146 57454
rect 240382 57218 249146 57454
rect 249382 57218 258146 57454
rect 258382 57218 267146 57454
rect 267382 57218 269708 57454
rect 269944 57218 270360 57454
rect 270596 57218 271166 57454
rect 271402 57218 280166 57454
rect 280402 57218 289166 57454
rect 289402 57218 298166 57454
rect 298402 57218 307166 57454
rect 307402 57218 309728 57454
rect 309964 57218 311380 57454
rect 311616 57218 312186 57454
rect 312422 57218 321186 57454
rect 321422 57218 330186 57454
rect 330422 57218 339186 57454
rect 339422 57218 348186 57454
rect 348422 57218 350748 57454
rect 350984 57218 352400 57454
rect 352636 57218 353206 57454
rect 353442 57218 362206 57454
rect 362442 57218 371206 57454
rect 371442 57218 380206 57454
rect 380442 57218 389206 57454
rect 389442 57218 391768 57454
rect 392004 57218 392420 57454
rect 392656 57218 393226 57454
rect 393462 57218 402226 57454
rect 402462 57218 411226 57454
rect 411462 57218 420226 57454
rect 420462 57218 429226 57454
rect 429462 57218 431788 57454
rect 432024 57218 432440 57454
rect 432676 57218 433246 57454
rect 433482 57218 442246 57454
rect 442482 57218 451246 57454
rect 451482 57218 460246 57454
rect 460482 57218 469246 57454
rect 469482 57218 471808 57454
rect 472044 57218 472460 57454
rect 472696 57218 473266 57454
rect 473502 57218 482266 57454
rect 482502 57218 491266 57454
rect 491502 57218 500266 57454
rect 500502 57218 509266 57454
rect 509502 57218 511828 57454
rect 512064 57218 512480 57454
rect 512716 57218 513286 57454
rect 513522 57218 522286 57454
rect 522522 57218 531286 57454
rect 531522 57218 540286 57454
rect 540522 57218 549286 57454
rect 549522 57218 551848 57454
rect 552084 57218 552500 57454
rect 552736 57218 553306 57454
rect 553542 57218 562306 57454
rect 562542 57218 571306 57454
rect 571542 57218 573836 57454
rect 574072 57218 579470 57454
rect 579706 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 4582 57134
rect 4818 56898 28240 57134
rect 28476 56898 29046 57134
rect 29282 56898 38046 57134
rect 38282 56898 47046 57134
rect 47282 56898 56046 57134
rect 56282 56898 65046 57134
rect 65282 56898 67608 57134
rect 67844 56898 68260 57134
rect 68496 56898 69066 57134
rect 69302 56898 78066 57134
rect 78302 56898 87066 57134
rect 87302 56898 96066 57134
rect 96302 56898 105066 57134
rect 105302 56898 107628 57134
rect 107864 56898 108280 57134
rect 108516 56898 109086 57134
rect 109322 56898 118086 57134
rect 118322 56898 127086 57134
rect 127322 56898 136086 57134
rect 136322 56898 145086 57134
rect 145322 56898 147648 57134
rect 147884 56898 149300 57134
rect 149536 56898 150106 57134
rect 150342 56898 159106 57134
rect 159342 56898 168106 57134
rect 168342 56898 177106 57134
rect 177342 56898 186106 57134
rect 186342 56898 188668 57134
rect 188904 56898 190320 57134
rect 190556 56898 191126 57134
rect 191362 56898 200126 57134
rect 200362 56898 209126 57134
rect 209362 56898 218126 57134
rect 218362 56898 227126 57134
rect 227362 56898 229688 57134
rect 229924 56898 230340 57134
rect 230576 56898 231146 57134
rect 231382 56898 240146 57134
rect 240382 56898 249146 57134
rect 249382 56898 258146 57134
rect 258382 56898 267146 57134
rect 267382 56898 269708 57134
rect 269944 56898 270360 57134
rect 270596 56898 271166 57134
rect 271402 56898 280166 57134
rect 280402 56898 289166 57134
rect 289402 56898 298166 57134
rect 298402 56898 307166 57134
rect 307402 56898 309728 57134
rect 309964 56898 311380 57134
rect 311616 56898 312186 57134
rect 312422 56898 321186 57134
rect 321422 56898 330186 57134
rect 330422 56898 339186 57134
rect 339422 56898 348186 57134
rect 348422 56898 350748 57134
rect 350984 56898 352400 57134
rect 352636 56898 353206 57134
rect 353442 56898 362206 57134
rect 362442 56898 371206 57134
rect 371442 56898 380206 57134
rect 380442 56898 389206 57134
rect 389442 56898 391768 57134
rect 392004 56898 392420 57134
rect 392656 56898 393226 57134
rect 393462 56898 402226 57134
rect 402462 56898 411226 57134
rect 411462 56898 420226 57134
rect 420462 56898 429226 57134
rect 429462 56898 431788 57134
rect 432024 56898 432440 57134
rect 432676 56898 433246 57134
rect 433482 56898 442246 57134
rect 442482 56898 451246 57134
rect 451482 56898 460246 57134
rect 460482 56898 469246 57134
rect 469482 56898 471808 57134
rect 472044 56898 472460 57134
rect 472696 56898 473266 57134
rect 473502 56898 482266 57134
rect 482502 56898 491266 57134
rect 491502 56898 500266 57134
rect 500502 56898 509266 57134
rect 509502 56898 511828 57134
rect 512064 56898 512480 57134
rect 512716 56898 513286 57134
rect 513522 56898 522286 57134
rect 522522 56898 531286 57134
rect 531522 56898 540286 57134
rect 540522 56898 549286 57134
rect 549522 56898 551848 57134
rect 552084 56898 552500 57134
rect 552736 56898 553306 57134
rect 553542 56898 562306 57134
rect 562542 56898 571306 57134
rect 571542 56898 573836 57134
rect 574072 56898 579470 57134
rect 579706 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 5382 39454
rect 5618 39218 578670 39454
rect 578906 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 5382 39134
rect 5618 38898 578670 39134
rect 578906 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use eFPGA_CPU_top  inst_eFPGA_CPU_top
timestamp 1637968891
transform 1 0 4000 0 1 30000
box 0 0 576288 648788
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 680788 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 680788 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 680788 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 680788 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 680788 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 680788 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 680788 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 680788 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 680788 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 680788 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 680788 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 680788 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 680788 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 680788 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 680788 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 680788 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 680788 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 680788 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 680788 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 680788 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 680788 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 680788 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 680788 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 680788 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 680788 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 680788 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 680788 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 680788 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 680788 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 680788 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 680788 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 680788 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 680788 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 680788 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 680788 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 680788 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 680788 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 680788 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 680788 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 680788 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 680788 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 680788 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 680788 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 680788 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 680788 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 680788 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 680788 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 680788 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 680788 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 680788 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 680788 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 680788 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 680788 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 680788 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 680788 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 680788 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 680788 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 680788 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 680788 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 680788 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 680788 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 680788 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 680788 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 680788 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 680788 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 680788 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 680788 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 680788 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 680788 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 680788 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 680788 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 680788 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 680788 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 680788 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 680788 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 680788 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 680788 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 680788 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 680788 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 680788 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 680788 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 680788 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 680788 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 680788 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 680788 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 680788 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 680788 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 680788 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 680788 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 680788 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 680788 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 680788 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 680788 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 680788 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 680788 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 680788 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 680788 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 680788 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 680788 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 680788 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 680788 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 680788 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 680788 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 680788 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 680788 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 680788 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 680788 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 680788 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 680788 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 680788 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 680788 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 680788 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 680788 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 680788 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 680788 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 680788 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 680788 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 680788 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 680788 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 680788 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 680788 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 680788 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 680788 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 680788 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 680788 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 680788 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 680788 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 680788 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 680788 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 680788 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
